module weight_lut (input logic clk, input logic [15:0] ind, output logic [15:0] out);

always_ff @ (negedge clk)
    case(ind)
    16'd0: out <= 16'hFFDA;    16'd1: out <= 16'hFB4B;    16'd2: out <= 16'hFCA5;    16'd3: out <= 16'h09A0;
    16'd4: out <= 16'hFE1B;    16'd5: out <= 16'h02FB;    16'd6: out <= 16'h01F1;    16'd7: out <= 16'h0264;
    16'd8: out <= 16'h0027;    16'd9: out <= 16'h0986;    16'd10: out <= 16'hFEA1;    16'd11: out <= 16'hF856;
    16'd12: out <= 16'h0078;    16'd13: out <= 16'hFA28;    16'd14: out <= 16'hFF21;    16'd15: out <= 16'hFB8B;
    16'd16: out <= 16'h010D;    16'd17: out <= 16'h050D;    16'd18: out <= 16'h0102;    16'd19: out <= 16'h0056;
    16'd20: out <= 16'h03C6;    16'd21: out <= 16'h026C;    16'd22: out <= 16'hFCFA;    16'd23: out <= 16'h01A9;
    16'd24: out <= 16'hFABB;    16'd25: out <= 16'h0358;    16'd26: out <= 16'h02D7;    16'd27: out <= 16'h01EB;
    16'd28: out <= 16'h0330;    16'd29: out <= 16'hFE7D;    16'd30: out <= 16'hFC20;    16'd31: out <= 16'hFE72;
    16'd32: out <= 16'h0517;    16'd33: out <= 16'hF925;    16'd34: out <= 16'hFFA4;    16'd35: out <= 16'h038D;
    16'd36: out <= 16'hFA8F;    16'd37: out <= 16'h0132;    16'd38: out <= 16'h007A;    16'd39: out <= 16'hFF33;
    16'd40: out <= 16'h0310;    16'd41: out <= 16'h015F;    16'd42: out <= 16'h0536;    16'd43: out <= 16'h008E;
    16'd44: out <= 16'hFDD6;    16'd45: out <= 16'hFD1C;    16'd46: out <= 16'hFA02;    16'd47: out <= 16'hFE00;
    16'd48: out <= 16'hFE3A;    16'd49: out <= 16'hFDA0;    16'd50: out <= 16'h055F;    16'd51: out <= 16'hFEAC;
    16'd52: out <= 16'h0525;    16'd53: out <= 16'hFED5;    16'd54: out <= 16'h0266;    16'd55: out <= 16'h070D;
    16'd56: out <= 16'hF784;    16'd57: out <= 16'h01BC;    16'd58: out <= 16'hFFDF;    16'd59: out <= 16'hFF7C;
    16'd60: out <= 16'h07FC;    16'd61: out <= 16'hF97C;    16'd62: out <= 16'hFF90;    16'd63: out <= 16'h0300;
    16'd64: out <= 16'hFF94;    16'd65: out <= 16'hFD50;    16'd66: out <= 16'h035C;    16'd67: out <= 16'h0244;
    16'd68: out <= 16'hF89B;    16'd69: out <= 16'hFF81;    16'd70: out <= 16'h0479;    16'd71: out <= 16'hFE75;
    16'd72: out <= 16'h03FA;    16'd73: out <= 16'h01A7;    16'd74: out <= 16'h01ED;    16'd75: out <= 16'hFFBE;
    16'd76: out <= 16'hFF18;    16'd77: out <= 16'h028B;    16'd78: out <= 16'hFBAC;    16'd79: out <= 16'hFCA7;
    16'd80: out <= 16'hFCFA;    16'd81: out <= 16'hFFCE;    16'd82: out <= 16'hFE68;    16'd83: out <= 16'hFDF0;
    16'd84: out <= 16'h0264;    16'd85: out <= 16'h0264;    16'd86: out <= 16'hF992;    16'd87: out <= 16'hFEBA;
    16'd88: out <= 16'h05BE;    16'd89: out <= 16'hFF82;    16'd90: out <= 16'h016D;    16'd91: out <= 16'h0345;
    16'd92: out <= 16'h0072;    16'd93: out <= 16'h011C;    16'd94: out <= 16'h0270;    16'd95: out <= 16'h01A0;
    16'd96: out <= 16'h0179;    16'd97: out <= 16'hFEDC;    16'd98: out <= 16'hFF57;    16'd99: out <= 16'h021B;
    16'd100: out <= 16'h004D;    16'd101: out <= 16'hFC21;    16'd102: out <= 16'h051C;    16'd103: out <= 16'hFE61;
    16'd104: out <= 16'hFE8B;    16'd105: out <= 16'h0185;    16'd106: out <= 16'h05AD;    16'd107: out <= 16'hFCF0;
    16'd108: out <= 16'hFEE4;    16'd109: out <= 16'hFFBD;    16'd110: out <= 16'hFA95;    16'd111: out <= 16'h0ACD;
    16'd112: out <= 16'hFC68;    16'd113: out <= 16'h002D;    16'd114: out <= 16'h038E;    16'd115: out <= 16'h0496;
    16'd116: out <= 16'hFC44;    16'd117: out <= 16'hFCDF;    16'd118: out <= 16'hFD54;    16'd119: out <= 16'hFFEC;
    16'd120: out <= 16'hFF68;    16'd121: out <= 16'h0592;    16'd122: out <= 16'hF725;    16'd123: out <= 16'h0379;
    16'd124: out <= 16'h06D5;    16'd125: out <= 16'h006A;    16'd126: out <= 16'hFE86;    16'd127: out <= 16'hFFE4;
    16'd128: out <= 16'h0370;    16'd129: out <= 16'h06B7;    16'd130: out <= 16'hFE0B;    16'd131: out <= 16'hFE9D;
    16'd132: out <= 16'hFD11;    16'd133: out <= 16'hFD50;    16'd134: out <= 16'hFF2B;    16'd135: out <= 16'hFD54;
    16'd136: out <= 16'h022E;    16'd137: out <= 16'h012C;    16'd138: out <= 16'hFFEB;    16'd139: out <= 16'hFB5B;
    16'd140: out <= 16'hFBF0;    16'd141: out <= 16'h048E;    16'd142: out <= 16'h020F;    16'd143: out <= 16'h03B9;
    16'd144: out <= 16'hFA45;    16'd145: out <= 16'h032E;    16'd146: out <= 16'h0596;    16'd147: out <= 16'h0300;
    16'd148: out <= 16'hFE4B;    16'd149: out <= 16'hFDB8;    16'd150: out <= 16'hFFFB;    16'd151: out <= 16'h01F3;
    16'd152: out <= 16'hFE35;    16'd153: out <= 16'h016A;    16'd154: out <= 16'hFD6A;    16'd155: out <= 16'hFD98;
    16'd156: out <= 16'hFD22;    16'd157: out <= 16'h0694;    16'd158: out <= 16'hFC53;    16'd159: out <= 16'hFE97;
    16'd160: out <= 16'hFAA9;    16'd161: out <= 16'hFD25;    16'd162: out <= 16'h02A1;    16'd163: out <= 16'hFA30;
    16'd164: out <= 16'h0326;    16'd165: out <= 16'h078E;    16'd166: out <= 16'h01F1;    16'd167: out <= 16'h01D3;
    16'd168: out <= 16'h028E;    16'd169: out <= 16'h09BE;    16'd170: out <= 16'h02BE;    16'd171: out <= 16'hFEEE;
    16'd172: out <= 16'hFDE3;    16'd173: out <= 16'h04E5;    16'd174: out <= 16'h043E;    16'd175: out <= 16'hFF5C;
    16'd176: out <= 16'hFF7C;    16'd177: out <= 16'hFF32;    16'd178: out <= 16'hFF16;    16'd179: out <= 16'hFF88;
    16'd180: out <= 16'hFE09;    16'd181: out <= 16'hFAB2;    16'd182: out <= 16'h0176;    16'd183: out <= 16'h055B;
    16'd184: out <= 16'h0861;    16'd185: out <= 16'hFA10;    16'd186: out <= 16'hFC93;    16'd187: out <= 16'h0060;
    16'd188: out <= 16'hFA21;    16'd189: out <= 16'hFFAE;    16'd190: out <= 16'h027F;    16'd191: out <= 16'hFCC0;
    16'd192: out <= 16'h0458;    16'd193: out <= 16'h085E;    16'd194: out <= 16'h0006;    16'd195: out <= 16'h008B;
    16'd196: out <= 16'h0235;    16'd197: out <= 16'hFD50;    16'd198: out <= 16'h03A4;    16'd199: out <= 16'hFE98;
    16'd200: out <= 16'h06DC;    16'd201: out <= 16'hFF2C;    16'd202: out <= 16'hFECC;    16'd203: out <= 16'hFF76;
    16'd204: out <= 16'hFFD9;    16'd205: out <= 16'h033A;    16'd206: out <= 16'h0502;    16'd207: out <= 16'h00A7;
    16'd208: out <= 16'hFC82;    16'd209: out <= 16'hFB15;    16'd210: out <= 16'hFE3A;    16'd211: out <= 16'hF9B5;
    16'd212: out <= 16'h03E2;    16'd213: out <= 16'hFC88;    16'd214: out <= 16'h02F9;    16'd215: out <= 16'hFF5B;
    16'd216: out <= 16'hFCCF;    16'd217: out <= 16'hFEF5;    16'd218: out <= 16'h004A;    16'd219: out <= 16'h0703;
    16'd220: out <= 16'hFE42;    16'd221: out <= 16'h0395;    16'd222: out <= 16'h0516;    16'd223: out <= 16'hFEAF;
    16'd224: out <= 16'hFBC2;    16'd225: out <= 16'hFD65;    16'd226: out <= 16'h0028;    16'd227: out <= 16'hFD7A;
    16'd228: out <= 16'hFFC9;    16'd229: out <= 16'h0261;    16'd230: out <= 16'hFE15;    16'd231: out <= 16'hF6EF;
    16'd232: out <= 16'h047D;    16'd233: out <= 16'hFAD0;    16'd234: out <= 16'h037B;    16'd235: out <= 16'hFDF8;
    16'd236: out <= 16'hFBDB;    16'd237: out <= 16'hFD26;    16'd238: out <= 16'h02D9;    16'd239: out <= 16'h0440;
    16'd240: out <= 16'hFFD4;    16'd241: out <= 16'hFFA5;    16'd242: out <= 16'hFC57;    16'd243: out <= 16'hFE1F;
    16'd244: out <= 16'hFD14;    16'd245: out <= 16'h031C;    16'd246: out <= 16'hFBBD;    16'd247: out <= 16'h062B;
    16'd248: out <= 16'h0123;    16'd249: out <= 16'h01BE;    16'd250: out <= 16'hFA73;    16'd251: out <= 16'h0A3C;
    16'd252: out <= 16'hF805;    16'd253: out <= 16'h0453;    16'd254: out <= 16'h0059;    16'd255: out <= 16'hFFEB;
    16'd256: out <= 16'hFAD5;    16'd257: out <= 16'h00FD;    16'd258: out <= 16'h0B5D;    16'd259: out <= 16'hFF19;
    16'd260: out <= 16'h02F9;    16'd261: out <= 16'hF952;    16'd262: out <= 16'hFD58;    16'd263: out <= 16'hF44C;
    16'd264: out <= 16'hFF22;    16'd265: out <= 16'hFF5C;    16'd266: out <= 16'h02D3;    16'd267: out <= 16'hFD19;
    16'd268: out <= 16'h064B;    16'd269: out <= 16'hFA74;    16'd270: out <= 16'hFF62;    16'd271: out <= 16'h01FE;
    16'd272: out <= 16'hFA7A;    16'd273: out <= 16'h016A;    16'd274: out <= 16'h00BA;    16'd275: out <= 16'h036B;
    16'd276: out <= 16'hFB42;    16'd277: out <= 16'h0278;    16'd278: out <= 16'hFF81;    16'd279: out <= 16'h05E4;
    16'd280: out <= 16'hFA1D;    16'd281: out <= 16'h06B4;    16'd282: out <= 16'h025A;    16'd283: out <= 16'hFEC3;
    16'd284: out <= 16'hFFF9;    16'd285: out <= 16'h01D0;    16'd286: out <= 16'h00F6;    16'd287: out <= 16'hFDAD;
    16'd288: out <= 16'h0473;    16'd289: out <= 16'hFF3E;    16'd290: out <= 16'h0482;    16'd291: out <= 16'h00B9;
    16'd292: out <= 16'h01D5;    16'd293: out <= 16'h0A15;    16'd294: out <= 16'h00B1;    16'd295: out <= 16'h05FE;
    16'd296: out <= 16'hFE1F;    16'd297: out <= 16'hFFE8;    16'd298: out <= 16'hFE94;    16'd299: out <= 16'hF8D2;
    16'd300: out <= 16'h03F1;    16'd301: out <= 16'h02E0;    16'd302: out <= 16'hFF51;    16'd303: out <= 16'h0012;
    16'd304: out <= 16'hFBC0;    16'd305: out <= 16'h0128;    16'd306: out <= 16'h010A;    16'd307: out <= 16'h06D0;
    16'd308: out <= 16'hFF3B;    16'd309: out <= 16'h03AF;    16'd310: out <= 16'h04D5;    16'd311: out <= 16'hFDCB;
    16'd312: out <= 16'hF71A;    16'd313: out <= 16'h0355;    16'd314: out <= 16'h044B;    16'd315: out <= 16'h0227;
    16'd316: out <= 16'hFF95;    16'd317: out <= 16'h013A;    16'd318: out <= 16'h0379;    16'd319: out <= 16'hFF0D;
    16'd320: out <= 16'hFC52;    16'd321: out <= 16'hFF42;    16'd322: out <= 16'h0362;    16'd323: out <= 16'h0423;
    16'd324: out <= 16'hFD8D;    16'd325: out <= 16'hFBD6;    16'd326: out <= 16'hFCB8;    16'd327: out <= 16'hFD4D;
    16'd328: out <= 16'hFE44;    16'd329: out <= 16'hFB8D;    16'd330: out <= 16'h0074;    16'd331: out <= 16'hFD7A;
    16'd332: out <= 16'h0091;    16'd333: out <= 16'hFFB9;    16'd334: out <= 16'hFCD9;    16'd335: out <= 16'hF99C;
    16'd336: out <= 16'h0059;    16'd337: out <= 16'hFC22;    16'd338: out <= 16'h00CD;    16'd339: out <= 16'hFECD;
    16'd340: out <= 16'hFAEE;    16'd341: out <= 16'h0406;    16'd342: out <= 16'hFD08;    16'd343: out <= 16'hFB33;
    16'd344: out <= 16'h053D;    16'd345: out <= 16'h0188;    16'd346: out <= 16'h033C;    16'd347: out <= 16'h03BF;
    16'd348: out <= 16'hFC33;    16'd349: out <= 16'h0188;    16'd350: out <= 16'h006F;    16'd351: out <= 16'h0045;
    16'd352: out <= 16'h051E;    16'd353: out <= 16'h00C3;    16'd354: out <= 16'hFCD7;    16'd355: out <= 16'h033F;
    16'd356: out <= 16'h02DE;    16'd357: out <= 16'hFA4E;    16'd358: out <= 16'hF41C;    16'd359: out <= 16'h01CD;
    16'd360: out <= 16'hFE37;    16'd361: out <= 16'hFDA0;    16'd362: out <= 16'hFECE;    16'd363: out <= 16'h04B1;
    16'd364: out <= 16'hFE40;    16'd365: out <= 16'h01AA;    16'd366: out <= 16'h01E9;    16'd367: out <= 16'hFECC;
    16'd368: out <= 16'h0481;    16'd369: out <= 16'h012F;    16'd370: out <= 16'h066D;    16'd371: out <= 16'h02EA;
    16'd372: out <= 16'hFFFD;    16'd373: out <= 16'hFF3E;    16'd374: out <= 16'hFD90;    16'd375: out <= 16'h05AA;
    16'd376: out <= 16'hFE29;    16'd377: out <= 16'hF6A3;    16'd378: out <= 16'hFDB7;    16'd379: out <= 16'hFDF1;
    16'd380: out <= 16'h0101;    16'd381: out <= 16'h094B;    16'd382: out <= 16'hFC66;    16'd383: out <= 16'h0450;
    16'd384: out <= 16'hFEEA;    16'd385: out <= 16'h0013;    16'd386: out <= 16'hFE35;    16'd387: out <= 16'hFF60;
    16'd388: out <= 16'h08CC;    16'd389: out <= 16'hFFE6;    16'd390: out <= 16'hFF89;    16'd391: out <= 16'h0085;
    16'd392: out <= 16'hFDD4;    16'd393: out <= 16'h00BB;    16'd394: out <= 16'hFE76;    16'd395: out <= 16'hFD99;
    16'd396: out <= 16'hFDC8;    16'd397: out <= 16'hFD9A;    16'd398: out <= 16'hFD04;    16'd399: out <= 16'h0036;
    16'd400: out <= 16'hFC95;    16'd401: out <= 16'h02F7;    16'd402: out <= 16'hFFB8;    16'd403: out <= 16'hFD0D;
    16'd404: out <= 16'hF858;    16'd405: out <= 16'h00A2;    16'd406: out <= 16'hFE40;    16'd407: out <= 16'hFDF2;
    16'd408: out <= 16'h02FD;    16'd409: out <= 16'h0807;    16'd410: out <= 16'h047F;    16'd411: out <= 16'h0244;
    16'd412: out <= 16'hFF75;    16'd413: out <= 16'hFFBE;    16'd414: out <= 16'hFBCB;    16'd415: out <= 16'hFE66;
    16'd416: out <= 16'hFFA4;    16'd417: out <= 16'hF90D;    16'd418: out <= 16'hFEE4;    16'd419: out <= 16'h016D;
    16'd420: out <= 16'h01A4;    16'd421: out <= 16'hFEF0;    16'd422: out <= 16'hF216;    16'd423: out <= 16'hFC57;
    16'd424: out <= 16'h0263;    16'd425: out <= 16'hFCA6;    16'd426: out <= 16'hFEAC;    16'd427: out <= 16'hFC30;
    16'd428: out <= 16'hFBFD;    16'd429: out <= 16'hFE8B;    16'd430: out <= 16'hFDEC;    16'd431: out <= 16'hF818;
    16'd432: out <= 16'h0221;    16'd433: out <= 16'hFE45;    16'd434: out <= 16'hFC62;    16'd435: out <= 16'hFA45;
    16'd436: out <= 16'hFE96;    16'd437: out <= 16'h031B;    16'd438: out <= 16'hFC82;    16'd439: out <= 16'h0513;
    16'd440: out <= 16'h044F;    16'd441: out <= 16'hFBC7;    16'd442: out <= 16'h021B;    16'd443: out <= 16'hFDD9;
    16'd444: out <= 16'hFD68;    16'd445: out <= 16'h0181;    16'd446: out <= 16'h0389;    16'd447: out <= 16'hFFDD;
    16'd448: out <= 16'hFEF9;    16'd449: out <= 16'hFF24;    16'd450: out <= 16'h0934;    16'd451: out <= 16'hFC62;
    16'd452: out <= 16'h0229;    16'd453: out <= 16'hFEC5;    16'd454: out <= 16'h04B2;    16'd455: out <= 16'hFE88;
    16'd456: out <= 16'h024E;    16'd457: out <= 16'h0288;    16'd458: out <= 16'h0037;    16'd459: out <= 16'hFC87;
    16'd460: out <= 16'hF9D4;    16'd461: out <= 16'hFE43;    16'd462: out <= 16'h09D3;    16'd463: out <= 16'hFE86;
    16'd464: out <= 16'hFDCB;    16'd465: out <= 16'h01D1;    16'd466: out <= 16'hF917;    16'd467: out <= 16'h03BD;
    16'd468: out <= 16'hFC5B;    16'd469: out <= 16'hFBD6;    16'd470: out <= 16'hF6A8;    16'd471: out <= 16'hFC7A;
    16'd472: out <= 16'hF80C;    16'd473: out <= 16'h00C0;    16'd474: out <= 16'h04CA;    16'd475: out <= 16'hFE97;
    16'd476: out <= 16'h0244;    16'd477: out <= 16'h055F;    16'd478: out <= 16'h00E7;    16'd479: out <= 16'hFDF7;
    16'd480: out <= 16'hFF4F;    16'd481: out <= 16'hF932;    16'd482: out <= 16'hFD0B;    16'd483: out <= 16'hFD5E;
    16'd484: out <= 16'h0573;    16'd485: out <= 16'hFB5E;    16'd486: out <= 16'hFDF1;    16'd487: out <= 16'hF9F2;
    16'd488: out <= 16'hF728;    16'd489: out <= 16'hFCA9;    16'd490: out <= 16'h02E7;    16'd491: out <= 16'hFEC9;
    16'd492: out <= 16'h0029;    16'd493: out <= 16'h0552;    16'd494: out <= 16'hFD6C;    16'd495: out <= 16'h00E0;
    16'd496: out <= 16'h0258;    16'd497: out <= 16'hFF2F;    16'd498: out <= 16'hFABE;    16'd499: out <= 16'h0348;
    16'd500: out <= 16'h0252;    16'd501: out <= 16'hFDE4;    16'd502: out <= 16'hFB13;    16'd503: out <= 16'hFC60;
    16'd504: out <= 16'hFC79;    16'd505: out <= 16'hFB4D;    16'd506: out <= 16'h012F;    16'd507: out <= 16'h03E5;
    16'd508: out <= 16'h022A;    16'd509: out <= 16'h0A22;    16'd510: out <= 16'hF997;    16'd511: out <= 16'h01B3;
    16'd512: out <= 16'h0210;    16'd513: out <= 16'hFBFF;    16'd514: out <= 16'h02F7;    16'd515: out <= 16'hFDDD;
    16'd516: out <= 16'h00FD;    16'd517: out <= 16'h0183;    16'd518: out <= 16'h0519;    16'd519: out <= 16'hFCBF;
    16'd520: out <= 16'h04D7;    16'd521: out <= 16'hF7D4;    16'd522: out <= 16'hFBAD;    16'd523: out <= 16'h0222;
    16'd524: out <= 16'hFC66;    16'd525: out <= 16'h0217;    16'd526: out <= 16'hFE4D;    16'd527: out <= 16'hF919;
    16'd528: out <= 16'hF6DD;    16'd529: out <= 16'h035E;    16'd530: out <= 16'h0D33;    16'd531: out <= 16'hFC99;
    16'd532: out <= 16'hFDC1;    16'd533: out <= 16'h06C6;    16'd534: out <= 16'h06FF;    16'd535: out <= 16'h0178;
    16'd536: out <= 16'h018B;    16'd537: out <= 16'hFC4D;    16'd538: out <= 16'h064A;    16'd539: out <= 16'hFEEE;
    16'd540: out <= 16'h0535;    16'd541: out <= 16'hFCD3;    16'd542: out <= 16'hFEF8;    16'd543: out <= 16'hFD63;
    16'd544: out <= 16'h02EB;    16'd545: out <= 16'hFCED;    16'd546: out <= 16'hFCB2;    16'd547: out <= 16'h0C9E;
    16'd548: out <= 16'h0470;    16'd549: out <= 16'hFAB5;    16'd550: out <= 16'h052E;    16'd551: out <= 16'hFE60;
    16'd552: out <= 16'hFE05;    16'd553: out <= 16'hFDAE;    16'd554: out <= 16'h060A;    16'd555: out <= 16'h006B;
    16'd556: out <= 16'h0409;    16'd557: out <= 16'h09A6;    16'd558: out <= 16'h00D9;    16'd559: out <= 16'hFE99;
    16'd560: out <= 16'h073B;    16'd561: out <= 16'hFAC2;    16'd562: out <= 16'h0266;    16'd563: out <= 16'h0047;
    16'd564: out <= 16'hFD0A;    16'd565: out <= 16'h0AB3;    16'd566: out <= 16'h0290;    16'd567: out <= 16'h00C2;
    16'd568: out <= 16'h0379;    16'd569: out <= 16'hFBBE;    16'd570: out <= 16'hFE07;    16'd571: out <= 16'h05F5;
    16'd572: out <= 16'hFE27;    16'd573: out <= 16'hF84B;    16'd574: out <= 16'h076B;    16'd575: out <= 16'h0359;
    16'd576: out <= 16'hFF9D;    16'd577: out <= 16'h0369;    16'd578: out <= 16'h01E1;    16'd579: out <= 16'h02E0;
    16'd580: out <= 16'h0293;    16'd581: out <= 16'hFE44;    16'd582: out <= 16'hFA53;    16'd583: out <= 16'h0140;
    16'd584: out <= 16'hFC53;    16'd585: out <= 16'h01C9;    16'd586: out <= 16'h06F7;    16'd587: out <= 16'hFCA9;
    16'd588: out <= 16'hFFC0;    16'd589: out <= 16'h0355;    16'd590: out <= 16'hFB59;    16'd591: out <= 16'h01A6;
    16'd592: out <= 16'h054D;    16'd593: out <= 16'hFF0B;    16'd594: out <= 16'h0149;    16'd595: out <= 16'hFE0C;
    16'd596: out <= 16'hFF6F;    16'd597: out <= 16'h0128;    16'd598: out <= 16'h0202;    16'd599: out <= 16'h0326;
    16'd600: out <= 16'hFDD2;    16'd601: out <= 16'h0483;    16'd602: out <= 16'hFD6C;    16'd603: out <= 16'hFC53;
    16'd604: out <= 16'h0247;    16'd605: out <= 16'h0297;    16'd606: out <= 16'hFCB4;    16'd607: out <= 16'hF92D;
    16'd608: out <= 16'h0996;    16'd609: out <= 16'hF813;    16'd610: out <= 16'h0173;    16'd611: out <= 16'h0209;
    16'd612: out <= 16'h0622;    16'd613: out <= 16'h0082;    16'd614: out <= 16'h014B;    16'd615: out <= 16'hFDFA;
    16'd616: out <= 16'hFD2D;    16'd617: out <= 16'hFAA8;    16'd618: out <= 16'h01B0;    16'd619: out <= 16'hFAEE;
    16'd620: out <= 16'h06E8;    16'd621: out <= 16'hFC1D;    16'd622: out <= 16'hFA7B;    16'd623: out <= 16'hFDEE;
    16'd624: out <= 16'hFE15;    16'd625: out <= 16'h023F;    16'd626: out <= 16'hFA6A;    16'd627: out <= 16'hF866;
    16'd628: out <= 16'hFAF5;    16'd629: out <= 16'h033C;    16'd630: out <= 16'h0853;    16'd631: out <= 16'h015C;
    16'd632: out <= 16'hFD81;    16'd633: out <= 16'hFE8D;    16'd634: out <= 16'h01CA;    16'd635: out <= 16'h00A9;
    16'd636: out <= 16'hFE9C;    16'd637: out <= 16'hFC47;    16'd638: out <= 16'hF3F1;    16'd639: out <= 16'h0017;
    16'd640: out <= 16'hFFA0;    16'd641: out <= 16'hFE9D;    16'd642: out <= 16'h05F8;    16'd643: out <= 16'h02EB;
    16'd644: out <= 16'h0385;    16'd645: out <= 16'hF7BE;    16'd646: out <= 16'h00B4;    16'd647: out <= 16'hFDEB;
    16'd648: out <= 16'hFA27;    16'd649: out <= 16'hFC82;    16'd650: out <= 16'hFB85;    16'd651: out <= 16'hFDD0;
    16'd652: out <= 16'hFF69;    16'd653: out <= 16'h03F9;    16'd654: out <= 16'h0407;    16'd655: out <= 16'hFAA1;
    16'd656: out <= 16'hFDA4;    16'd657: out <= 16'hFD63;    16'd658: out <= 16'h0096;    16'd659: out <= 16'hFF01;
    16'd660: out <= 16'hF912;    16'd661: out <= 16'hFC92;    16'd662: out <= 16'h01B9;    16'd663: out <= 16'hFB30;
    16'd664: out <= 16'h0210;    16'd665: out <= 16'hFA74;    16'd666: out <= 16'hFAD0;    16'd667: out <= 16'hFFB5;
    16'd668: out <= 16'hFEAD;    16'd669: out <= 16'h00A8;    16'd670: out <= 16'hFAB0;    16'd671: out <= 16'hFA7D;
    16'd672: out <= 16'h07F4;    16'd673: out <= 16'hFE00;    16'd674: out <= 16'hF31D;    16'd675: out <= 16'hFE1A;
    16'd676: out <= 16'h02E6;    16'd677: out <= 16'h032C;    16'd678: out <= 16'hFC67;    16'd679: out <= 16'h028E;
    16'd680: out <= 16'h00C5;    16'd681: out <= 16'h017D;    16'd682: out <= 16'hFD12;    16'd683: out <= 16'hFA7E;
    16'd684: out <= 16'h0416;    16'd685: out <= 16'h0558;    16'd686: out <= 16'h032C;    16'd687: out <= 16'hFD1F;
    16'd688: out <= 16'hF945;    16'd689: out <= 16'h0199;    16'd690: out <= 16'hFFC1;    16'd691: out <= 16'hFFC7;
    16'd692: out <= 16'hFE85;    16'd693: out <= 16'hFF95;    16'd694: out <= 16'hFC72;    16'd695: out <= 16'h013C;
    16'd696: out <= 16'hFE0D;    16'd697: out <= 16'h085A;    16'd698: out <= 16'h0026;    16'd699: out <= 16'hFDBA;
    16'd700: out <= 16'hFD3F;    16'd701: out <= 16'h05D4;    16'd702: out <= 16'hFF3B;    16'd703: out <= 16'hFC38;
    16'd704: out <= 16'hFBFA;    16'd705: out <= 16'h04AF;    16'd706: out <= 16'h0488;    16'd707: out <= 16'hFDC4;
    16'd708: out <= 16'hFF4C;    16'd709: out <= 16'h037D;    16'd710: out <= 16'hF8C5;    16'd711: out <= 16'hFECD;
    16'd712: out <= 16'h02C3;    16'd713: out <= 16'hF863;    16'd714: out <= 16'h0258;    16'd715: out <= 16'h027B;
    16'd716: out <= 16'hFD57;    16'd717: out <= 16'hFE8B;    16'd718: out <= 16'h009F;    16'd719: out <= 16'hFEC3;
    16'd720: out <= 16'hFDE0;    16'd721: out <= 16'hF903;    16'd722: out <= 16'hF84F;    16'd723: out <= 16'hFD58;
    16'd724: out <= 16'hFE63;    16'd725: out <= 16'h01CF;    16'd726: out <= 16'h048C;    16'd727: out <= 16'h035E;
    16'd728: out <= 16'h0361;    16'd729: out <= 16'h003E;    16'd730: out <= 16'hFAF5;    16'd731: out <= 16'h06AB;
    16'd732: out <= 16'h05C0;    16'd733: out <= 16'hFD46;    16'd734: out <= 16'hFD22;    16'd735: out <= 16'hFD7B;
    16'd736: out <= 16'hFE75;    16'd737: out <= 16'h05C2;    16'd738: out <= 16'hFBA7;    16'd739: out <= 16'h0265;
    16'd740: out <= 16'hFDD9;    16'd741: out <= 16'h0456;    16'd742: out <= 16'hFE6F;    16'd743: out <= 16'hFD7A;
    16'd744: out <= 16'hFE97;    16'd745: out <= 16'hFDCD;    16'd746: out <= 16'hF8D8;    16'd747: out <= 16'hFF69;
    16'd748: out <= 16'hFD56;    16'd749: out <= 16'h00BE;    16'd750: out <= 16'h05BE;    16'd751: out <= 16'hFE5D;
    16'd752: out <= 16'hFBF0;    16'd753: out <= 16'h0495;    16'd754: out <= 16'hFD8D;    16'd755: out <= 16'h04BE;
    16'd756: out <= 16'hFB14;    16'd757: out <= 16'hFCF5;    16'd758: out <= 16'hFCF8;    16'd759: out <= 16'hFD29;
    16'd760: out <= 16'hFDBC;    16'd761: out <= 16'h04CE;    16'd762: out <= 16'hF694;    16'd763: out <= 16'hF9D3;
    16'd764: out <= 16'h011D;    16'd765: out <= 16'hFD21;    16'd766: out <= 16'hFE0A;    16'd767: out <= 16'h0111;
    16'd768: out <= 16'h05D2;    16'd769: out <= 16'hFD4B;    16'd770: out <= 16'hFD69;    16'd771: out <= 16'hFF72;
    16'd772: out <= 16'h030B;    16'd773: out <= 16'h0202;    16'd774: out <= 16'h02B5;    16'd775: out <= 16'h0270;
    16'd776: out <= 16'h01A6;    16'd777: out <= 16'hFA30;    16'd778: out <= 16'h0186;    16'd779: out <= 16'h0302;
    16'd780: out <= 16'hFE74;    16'd781: out <= 16'h024E;    16'd782: out <= 16'hFC99;    16'd783: out <= 16'h02A2;
    16'd784: out <= 16'hFD4B;    16'd785: out <= 16'hFBA6;    16'd786: out <= 16'hFEB2;    16'd787: out <= 16'hFFD1;
    16'd788: out <= 16'hFD96;    16'd789: out <= 16'hFDAA;    16'd790: out <= 16'hFB4D;    16'd791: out <= 16'hFE11;
    16'd792: out <= 16'hFD69;    16'd793: out <= 16'h0273;    16'd794: out <= 16'h02C9;    16'd795: out <= 16'h01B1;
    16'd796: out <= 16'h03F3;    16'd797: out <= 16'h079B;    16'd798: out <= 16'h01C1;    16'd799: out <= 16'hFDB8;
    16'd800: out <= 16'h0508;    16'd801: out <= 16'h03E8;    16'd802: out <= 16'h04EB;    16'd803: out <= 16'hFC09;
    16'd804: out <= 16'hFD19;    16'd805: out <= 16'hFBD4;    16'd806: out <= 16'h04F1;    16'd807: out <= 16'h0598;
    16'd808: out <= 16'hFBBA;    16'd809: out <= 16'hFFE8;    16'd810: out <= 16'hFEBB;    16'd811: out <= 16'h00FC;
    16'd812: out <= 16'h0303;    16'd813: out <= 16'hFCBF;    16'd814: out <= 16'h01BF;    16'd815: out <= 16'hF758;
    16'd816: out <= 16'hFD92;    16'd817: out <= 16'h0161;    16'd818: out <= 16'hFD99;    16'd819: out <= 16'h01DB;
    16'd820: out <= 16'h0109;    16'd821: out <= 16'hFDB4;    16'd822: out <= 16'h0090;    16'd823: out <= 16'hFADD;
    16'd824: out <= 16'hFCE2;    16'd825: out <= 16'h02A1;    16'd826: out <= 16'hFE65;    16'd827: out <= 16'h016C;
    16'd828: out <= 16'h0058;    16'd829: out <= 16'hFCB1;    16'd830: out <= 16'hFDB0;    16'd831: out <= 16'h022A;
    16'd832: out <= 16'hFBC0;    16'd833: out <= 16'h0169;    16'd834: out <= 16'h0724;    16'd835: out <= 16'hFE70;
    16'd836: out <= 16'hFC70;    16'd837: out <= 16'hFF47;    16'd838: out <= 16'hFED5;    16'd839: out <= 16'h0023;
    16'd840: out <= 16'hFB8C;    16'd841: out <= 16'h012A;    16'd842: out <= 16'h030E;    16'd843: out <= 16'hFEB2;
    16'd844: out <= 16'h038A;    16'd845: out <= 16'hFC73;    16'd846: out <= 16'hFEDE;    16'd847: out <= 16'hFFD9;
    16'd848: out <= 16'hFDFD;    16'd849: out <= 16'hFF32;    16'd850: out <= 16'h010C;    16'd851: out <= 16'hFB6B;
    16'd852: out <= 16'h00C0;    16'd853: out <= 16'h0088;    16'd854: out <= 16'h068A;    16'd855: out <= 16'hFF40;
    16'd856: out <= 16'hFC48;    16'd857: out <= 16'h0A30;    16'd858: out <= 16'hFB84;    16'd859: out <= 16'hFD99;
    16'd860: out <= 16'h0301;    16'd861: out <= 16'h0113;    16'd862: out <= 16'hFEDB;    16'd863: out <= 16'h0092;
    16'd864: out <= 16'hFB60;    16'd865: out <= 16'hFFB6;    16'd866: out <= 16'h0175;    16'd867: out <= 16'h00C8;
    16'd868: out <= 16'hFEBB;    16'd869: out <= 16'h03A8;    16'd870: out <= 16'hFCD0;    16'd871: out <= 16'h0457;
    16'd872: out <= 16'hFE5B;    16'd873: out <= 16'hFAF9;    16'd874: out <= 16'hFA84;    16'd875: out <= 16'hFDE0;
    16'd876: out <= 16'h00C7;    16'd877: out <= 16'hFD9D;    16'd878: out <= 16'h0047;    16'd879: out <= 16'hFAD5;
    16'd880: out <= 16'h01F0;    16'd881: out <= 16'h004C;    16'd882: out <= 16'h0421;    16'd883: out <= 16'hFF52;
    16'd884: out <= 16'h029A;    16'd885: out <= 16'hFC81;    16'd886: out <= 16'h0115;    16'd887: out <= 16'hFE40;
    16'd888: out <= 16'hFC44;    16'd889: out <= 16'h0395;    16'd890: out <= 16'hFC1F;    16'd891: out <= 16'hFE23;
    16'd892: out <= 16'hFCFB;    16'd893: out <= 16'h03CB;    16'd894: out <= 16'hFF4B;    16'd895: out <= 16'hFCFA;
    16'd896: out <= 16'h00DC;    16'd897: out <= 16'hFE39;    16'd898: out <= 16'hFE5D;    16'd899: out <= 16'hF83E;
    16'd900: out <= 16'hFD89;    16'd901: out <= 16'h028D;    16'd902: out <= 16'h0223;    16'd903: out <= 16'h04B5;
    16'd904: out <= 16'hFF59;    16'd905: out <= 16'h03AF;    16'd906: out <= 16'h01D3;    16'd907: out <= 16'hFDF8;
    16'd908: out <= 16'h07CA;    16'd909: out <= 16'hFAF4;    16'd910: out <= 16'hFA0D;    16'd911: out <= 16'hFC79;
    16'd912: out <= 16'h006F;    16'd913: out <= 16'hFED6;    16'd914: out <= 16'hFE95;    16'd915: out <= 16'h0072;
    16'd916: out <= 16'hFE5D;    16'd917: out <= 16'h02D3;    16'd918: out <= 16'hFD3C;    16'd919: out <= 16'hFA4B;
    16'd920: out <= 16'h02CF;    16'd921: out <= 16'h0193;    16'd922: out <= 16'h034A;    16'd923: out <= 16'hFDAC;
    16'd924: out <= 16'h035B;    16'd925: out <= 16'hFA0F;    16'd926: out <= 16'hF91F;    16'd927: out <= 16'hFC8B;
    16'd928: out <= 16'hFC0D;    16'd929: out <= 16'h00D3;    16'd930: out <= 16'h02AC;    16'd931: out <= 16'hF9E2;
    16'd932: out <= 16'hFFC5;    16'd933: out <= 16'hFD31;    16'd934: out <= 16'hFB72;    16'd935: out <= 16'h00F7;
    16'd936: out <= 16'hFD78;    16'd937: out <= 16'hFF15;    16'd938: out <= 16'h023E;    16'd939: out <= 16'h0237;
    16'd940: out <= 16'h06EA;    16'd941: out <= 16'hFE00;    16'd942: out <= 16'hFF55;    16'd943: out <= 16'h03F6;
    16'd944: out <= 16'h0546;    16'd945: out <= 16'h094F;    16'd946: out <= 16'h08E3;    16'd947: out <= 16'hFCF4;
    16'd948: out <= 16'h05B4;    16'd949: out <= 16'hFE5E;    16'd950: out <= 16'h046D;    16'd951: out <= 16'h0305;
    16'd952: out <= 16'h01E2;    16'd953: out <= 16'hFF5F;    16'd954: out <= 16'h0227;    16'd955: out <= 16'hFF5D;
    16'd956: out <= 16'h01CB;    16'd957: out <= 16'hFEF7;    16'd958: out <= 16'hFEF1;    16'd959: out <= 16'h04AA;
    16'd960: out <= 16'h01BB;    16'd961: out <= 16'h0071;    16'd962: out <= 16'h021E;    16'd963: out <= 16'hFD71;
    16'd964: out <= 16'hF836;    16'd965: out <= 16'h00AB;    16'd966: out <= 16'h035C;    16'd967: out <= 16'hFF1D;
    16'd968: out <= 16'h02B7;    16'd969: out <= 16'h0072;    16'd970: out <= 16'h0B2B;    16'd971: out <= 16'hF921;
    16'd972: out <= 16'h016A;    16'd973: out <= 16'hFCFD;    16'd974: out <= 16'hFAA4;    16'd975: out <= 16'h012A;
    16'd976: out <= 16'h05F7;    16'd977: out <= 16'h02A6;    16'd978: out <= 16'h02B8;    16'd979: out <= 16'h01B6;
    16'd980: out <= 16'h05B7;    16'd981: out <= 16'h00E2;    16'd982: out <= 16'h015D;    16'd983: out <= 16'hFA53;
    16'd984: out <= 16'hFF94;    16'd985: out <= 16'h04DD;    16'd986: out <= 16'h0275;    16'd987: out <= 16'hFC77;
    16'd988: out <= 16'h05FF;    16'd989: out <= 16'hFFB2;    16'd990: out <= 16'h0173;    16'd991: out <= 16'h07F0;
    16'd992: out <= 16'hFFFA;    16'd993: out <= 16'h02E9;    16'd994: out <= 16'h0672;    16'd995: out <= 16'h0144;
    16'd996: out <= 16'h046C;    16'd997: out <= 16'h0514;    16'd998: out <= 16'h0606;    16'd999: out <= 16'h021C;
    16'd1000: out <= 16'hFE6A;    16'd1001: out <= 16'h04F8;    16'd1002: out <= 16'hFC8A;    16'd1003: out <= 16'h057D;
    16'd1004: out <= 16'h0208;    16'd1005: out <= 16'hFF57;    16'd1006: out <= 16'h068B;    16'd1007: out <= 16'hFD9C;
    16'd1008: out <= 16'hF9F6;    16'd1009: out <= 16'hFF36;    16'd1010: out <= 16'h0688;    16'd1011: out <= 16'hFE10;
    16'd1012: out <= 16'hFB07;    16'd1013: out <= 16'h06C2;    16'd1014: out <= 16'h0416;    16'd1015: out <= 16'h0572;
    16'd1016: out <= 16'h0146;    16'd1017: out <= 16'h05FF;    16'd1018: out <= 16'hFC20;    16'd1019: out <= 16'hFF9C;
    16'd1020: out <= 16'hFEE4;    16'd1021: out <= 16'hFAE1;    16'd1022: out <= 16'h047A;    16'd1023: out <= 16'hFFF9;
    16'd1024: out <= 16'hFF18;    16'd1025: out <= 16'hFDBA;    16'd1026: out <= 16'h0538;    16'd1027: out <= 16'h0013;
    16'd1028: out <= 16'hFC3A;    16'd1029: out <= 16'h0319;    16'd1030: out <= 16'hFE83;    16'd1031: out <= 16'h0561;
    16'd1032: out <= 16'hFFD8;    16'd1033: out <= 16'hFE1B;    16'd1034: out <= 16'h013E;    16'd1035: out <= 16'h05F7;
    16'd1036: out <= 16'hFC85;    16'd1037: out <= 16'h017F;    16'd1038: out <= 16'hFDD7;    16'd1039: out <= 16'hFFE5;
    16'd1040: out <= 16'h007F;    16'd1041: out <= 16'hFBA9;    16'd1042: out <= 16'h00C9;    16'd1043: out <= 16'hFCFB;
    16'd1044: out <= 16'hFA58;    16'd1045: out <= 16'hFCCD;    16'd1046: out <= 16'h0AC4;    16'd1047: out <= 16'hFF92;
    16'd1048: out <= 16'h0298;    16'd1049: out <= 16'hFFC5;    16'd1050: out <= 16'h0256;    16'd1051: out <= 16'h0916;
    16'd1052: out <= 16'hFDD0;    16'd1053: out <= 16'hFED4;    16'd1054: out <= 16'hFE7D;    16'd1055: out <= 16'hFDF8;
    16'd1056: out <= 16'h0476;    16'd1057: out <= 16'hFBB1;    16'd1058: out <= 16'hFD34;    16'd1059: out <= 16'hFFE3;
    16'd1060: out <= 16'h0460;    16'd1061: out <= 16'hFE54;    16'd1062: out <= 16'hFABA;    16'd1063: out <= 16'hFE38;
    16'd1064: out <= 16'hFEED;    16'd1065: out <= 16'hFC4E;    16'd1066: out <= 16'hFFB5;    16'd1067: out <= 16'hFCD5;
    16'd1068: out <= 16'hFB44;    16'd1069: out <= 16'h015B;    16'd1070: out <= 16'h028E;    16'd1071: out <= 16'h02A8;
    16'd1072: out <= 16'h0369;    16'd1073: out <= 16'h040E;    16'd1074: out <= 16'h0086;    16'd1075: out <= 16'hFF42;
    16'd1076: out <= 16'hF972;    16'd1077: out <= 16'hFD68;    16'd1078: out <= 16'hFCF1;    16'd1079: out <= 16'h004C;
    16'd1080: out <= 16'hFD90;    16'd1081: out <= 16'h03AB;    16'd1082: out <= 16'hFB5B;    16'd1083: out <= 16'h06B6;
    16'd1084: out <= 16'hFFEB;    16'd1085: out <= 16'hF9EC;    16'd1086: out <= 16'hFB62;    16'd1087: out <= 16'hFEED;
    16'd1088: out <= 16'hFD28;    16'd1089: out <= 16'h0068;    16'd1090: out <= 16'hFC66;    16'd1091: out <= 16'hF772;
    16'd1092: out <= 16'h03C2;    16'd1093: out <= 16'hFCB2;    16'd1094: out <= 16'h029A;    16'd1095: out <= 16'h0A1A;
    16'd1096: out <= 16'h047C;    16'd1097: out <= 16'h04BE;    16'd1098: out <= 16'hFFFA;    16'd1099: out <= 16'hFCFD;
    16'd1100: out <= 16'h00A5;    16'd1101: out <= 16'hF9DB;    16'd1102: out <= 16'h0508;    16'd1103: out <= 16'h00BA;
    16'd1104: out <= 16'hFF9C;    16'd1105: out <= 16'hFCBA;    16'd1106: out <= 16'h00E6;    16'd1107: out <= 16'h0508;
    16'd1108: out <= 16'hFB95;    16'd1109: out <= 16'h0A8E;    16'd1110: out <= 16'hFF34;    16'd1111: out <= 16'hFD3A;
    16'd1112: out <= 16'hFD17;    16'd1113: out <= 16'hFF17;    16'd1114: out <= 16'hFC65;    16'd1115: out <= 16'hFD98;
    16'd1116: out <= 16'h0793;    16'd1117: out <= 16'hFDC4;    16'd1118: out <= 16'h00A2;    16'd1119: out <= 16'h0819;
    16'd1120: out <= 16'h0593;    16'd1121: out <= 16'h0016;    16'd1122: out <= 16'h050E;    16'd1123: out <= 16'h09A1;
    16'd1124: out <= 16'hFFE7;    16'd1125: out <= 16'hFE8B;    16'd1126: out <= 16'hFDF2;    16'd1127: out <= 16'h007B;
    16'd1128: out <= 16'h0043;    16'd1129: out <= 16'hFF8C;    16'd1130: out <= 16'h03A8;    16'd1131: out <= 16'hFCCB;
    16'd1132: out <= 16'h00C9;    16'd1133: out <= 16'hFD99;    16'd1134: out <= 16'h0169;    16'd1135: out <= 16'h0073;
    16'd1136: out <= 16'hFA53;    16'd1137: out <= 16'hFE05;    16'd1138: out <= 16'hFE9E;    16'd1139: out <= 16'hFF51;
    16'd1140: out <= 16'hF926;    16'd1141: out <= 16'hFABD;    16'd1142: out <= 16'hFF46;    16'd1143: out <= 16'hFB3F;
    16'd1144: out <= 16'h0386;    16'd1145: out <= 16'hFDF3;    16'd1146: out <= 16'h01C9;    16'd1147: out <= 16'hFEC3;
    16'd1148: out <= 16'hFB22;    16'd1149: out <= 16'hF8BE;    16'd1150: out <= 16'h0148;    16'd1151: out <= 16'h0675;
    16'd1152: out <= 16'hFE71;    16'd1153: out <= 16'hFE61;    16'd1154: out <= 16'h0831;    16'd1155: out <= 16'h04C5;
    16'd1156: out <= 16'hFCC7;    16'd1157: out <= 16'hF539;    16'd1158: out <= 16'h0764;    16'd1159: out <= 16'h06BA;
    16'd1160: out <= 16'h01DD;    16'd1161: out <= 16'h0129;    16'd1162: out <= 16'h01C3;    16'd1163: out <= 16'hFB0F;
    16'd1164: out <= 16'hFD63;    16'd1165: out <= 16'h08B7;    16'd1166: out <= 16'hFD76;    16'd1167: out <= 16'hFC23;
    16'd1168: out <= 16'hFCA7;    16'd1169: out <= 16'hFE00;    16'd1170: out <= 16'hFAA3;    16'd1171: out <= 16'hFF65;
    16'd1172: out <= 16'h039D;    16'd1173: out <= 16'hFEFD;    16'd1174: out <= 16'h03D5;    16'd1175: out <= 16'hFF4F;
    16'd1176: out <= 16'h02A4;    16'd1177: out <= 16'hFAFC;    16'd1178: out <= 16'h02EC;    16'd1179: out <= 16'h0332;
    16'd1180: out <= 16'hFDEE;    16'd1181: out <= 16'hFE40;    16'd1182: out <= 16'h035B;    16'd1183: out <= 16'h06EE;
    16'd1184: out <= 16'h03ED;    16'd1185: out <= 16'h04F2;    16'd1186: out <= 16'h0437;    16'd1187: out <= 16'h02D0;
    16'd1188: out <= 16'hFA87;    16'd1189: out <= 16'hF407;    16'd1190: out <= 16'hFB12;    16'd1191: out <= 16'h0467;
    16'd1192: out <= 16'h04CA;    16'd1193: out <= 16'h02ED;    16'd1194: out <= 16'h07C5;    16'd1195: out <= 16'h0258;
    16'd1196: out <= 16'hFA23;    16'd1197: out <= 16'hF9FC;    16'd1198: out <= 16'h015E;    16'd1199: out <= 16'h00B3;
    16'd1200: out <= 16'hF5C8;    16'd1201: out <= 16'h02C0;    16'd1202: out <= 16'hFDCD;    16'd1203: out <= 16'hFE3A;
    16'd1204: out <= 16'h04E6;    16'd1205: out <= 16'hFFDA;    16'd1206: out <= 16'h0123;    16'd1207: out <= 16'h0328;
    16'd1208: out <= 16'h03DE;    16'd1209: out <= 16'h00F7;    16'd1210: out <= 16'h05FB;    16'd1211: out <= 16'hFD74;
    16'd1212: out <= 16'h010F;    16'd1213: out <= 16'hFCDE;    16'd1214: out <= 16'h0369;    16'd1215: out <= 16'hFD7D;
    16'd1216: out <= 16'hFBDD;    16'd1217: out <= 16'hFE04;    16'd1218: out <= 16'hF649;    16'd1219: out <= 16'hFE74;
    16'd1220: out <= 16'hFF87;    16'd1221: out <= 16'hF993;    16'd1222: out <= 16'h055C;    16'd1223: out <= 16'hFF11;
    16'd1224: out <= 16'hFF2D;    16'd1225: out <= 16'h0582;    16'd1226: out <= 16'h00CD;    16'd1227: out <= 16'hFD76;
    16'd1228: out <= 16'hFFEE;    16'd1229: out <= 16'h01E1;    16'd1230: out <= 16'hFB3E;    16'd1231: out <= 16'hFF32;
    16'd1232: out <= 16'hF95E;    16'd1233: out <= 16'hFF84;    16'd1234: out <= 16'h00EB;    16'd1235: out <= 16'h0352;
    16'd1236: out <= 16'hF92D;    16'd1237: out <= 16'h03B7;    16'd1238: out <= 16'hFFE3;    16'd1239: out <= 16'h03BF;
    16'd1240: out <= 16'hFCEE;    16'd1241: out <= 16'hFF59;    16'd1242: out <= 16'h03D0;    16'd1243: out <= 16'hFEBB;
    16'd1244: out <= 16'hFA0D;    16'd1245: out <= 16'h0148;    16'd1246: out <= 16'h02EA;    16'd1247: out <= 16'h0350;
    16'd1248: out <= 16'h062F;    16'd1249: out <= 16'hFE0D;    16'd1250: out <= 16'hFA7B;    16'd1251: out <= 16'h0392;
    16'd1252: out <= 16'h0330;    16'd1253: out <= 16'hFF0F;    16'd1254: out <= 16'hFF0E;    16'd1255: out <= 16'hFDFB;
    16'd1256: out <= 16'hFEA0;    16'd1257: out <= 16'hFAA4;    16'd1258: out <= 16'hFC09;    16'd1259: out <= 16'hFE14;
    16'd1260: out <= 16'hFF8F;    16'd1261: out <= 16'h068D;    16'd1262: out <= 16'hFE4E;    16'd1263: out <= 16'h00BD;
    16'd1264: out <= 16'hFF24;    16'd1265: out <= 16'hFBD1;    16'd1266: out <= 16'h00AD;    16'd1267: out <= 16'h00F5;
    16'd1268: out <= 16'h011D;    16'd1269: out <= 16'h097F;    16'd1270: out <= 16'h0230;    16'd1271: out <= 16'hFB51;
    16'd1272: out <= 16'h037C;    16'd1273: out <= 16'hFD51;    16'd1274: out <= 16'h0679;    16'd1275: out <= 16'h0000;
    16'd1276: out <= 16'h00EE;    16'd1277: out <= 16'h0082;    16'd1278: out <= 16'h082B;    16'd1279: out <= 16'hFE51;
    16'd1280: out <= 16'hFE66;    16'd1281: out <= 16'hFA5F;    16'd1282: out <= 16'hFC83;    16'd1283: out <= 16'h00FD;
    16'd1284: out <= 16'hFFE4;    16'd1285: out <= 16'hF7C3;    16'd1286: out <= 16'h03FA;    16'd1287: out <= 16'h0604;
    16'd1288: out <= 16'h00EC;    16'd1289: out <= 16'hF75E;    16'd1290: out <= 16'hFFF2;    16'd1291: out <= 16'hFF8E;
    16'd1292: out <= 16'hFFAB;    16'd1293: out <= 16'hFB44;    16'd1294: out <= 16'h0219;    16'd1295: out <= 16'h0235;
    16'd1296: out <= 16'hF7C1;    16'd1297: out <= 16'hFDD5;    16'd1298: out <= 16'hFB5C;    16'd1299: out <= 16'h0470;
    16'd1300: out <= 16'h027F;    16'd1301: out <= 16'h0295;    16'd1302: out <= 16'h04A8;    16'd1303: out <= 16'hFBA5;
    16'd1304: out <= 16'hFDD4;    16'd1305: out <= 16'h038B;    16'd1306: out <= 16'h03AD;    16'd1307: out <= 16'hFFEA;
    16'd1308: out <= 16'hFE44;    16'd1309: out <= 16'h034A;    16'd1310: out <= 16'h0332;    16'd1311: out <= 16'h06EF;
    16'd1312: out <= 16'hFF67;    16'd1313: out <= 16'hFE70;    16'd1314: out <= 16'hFBD6;    16'd1315: out <= 16'h016D;
    16'd1316: out <= 16'hFEBF;    16'd1317: out <= 16'hFEFF;    16'd1318: out <= 16'h0121;    16'd1319: out <= 16'h05CE;
    16'd1320: out <= 16'hFF5D;    16'd1321: out <= 16'h0006;    16'd1322: out <= 16'h0064;    16'd1323: out <= 16'h0543;
    16'd1324: out <= 16'h02E9;    16'd1325: out <= 16'hFD68;    16'd1326: out <= 16'hFB2F;    16'd1327: out <= 16'hFBC9;
    16'd1328: out <= 16'hFC32;    16'd1329: out <= 16'h0060;    16'd1330: out <= 16'hFC5B;    16'd1331: out <= 16'h0036;
    16'd1332: out <= 16'hFB00;    16'd1333: out <= 16'hFDFE;    16'd1334: out <= 16'hFBED;    16'd1335: out <= 16'h042A;
    16'd1336: out <= 16'hFDA5;    16'd1337: out <= 16'h00C2;    16'd1338: out <= 16'h0277;    16'd1339: out <= 16'h0871;
    16'd1340: out <= 16'h044D;    16'd1341: out <= 16'h006F;    16'd1342: out <= 16'h00CC;    16'd1343: out <= 16'h01AF;
    16'd1344: out <= 16'h0372;    16'd1345: out <= 16'hFD66;    16'd1346: out <= 16'hFE37;    16'd1347: out <= 16'h016E;
    16'd1348: out <= 16'hFD7A;    16'd1349: out <= 16'h0090;    16'd1350: out <= 16'h03AC;    16'd1351: out <= 16'hFD1F;
    16'd1352: out <= 16'h0258;    16'd1353: out <= 16'h024D;    16'd1354: out <= 16'hFF7F;    16'd1355: out <= 16'h0291;
    16'd1356: out <= 16'hFCFD;    16'd1357: out <= 16'h04B5;    16'd1358: out <= 16'hFEFD;    16'd1359: out <= 16'hFF81;
    16'd1360: out <= 16'h0380;    16'd1361: out <= 16'h0223;    16'd1362: out <= 16'h03B6;    16'd1363: out <= 16'h08F1;
    16'd1364: out <= 16'hFEF5;    16'd1365: out <= 16'h03BB;    16'd1366: out <= 16'h02AA;    16'd1367: out <= 16'hFFCD;
    16'd1368: out <= 16'h00EA;    16'd1369: out <= 16'h0088;    16'd1370: out <= 16'h0265;    16'd1371: out <= 16'hFE30;
    16'd1372: out <= 16'h02C3;    16'd1373: out <= 16'h0582;    16'd1374: out <= 16'hFB73;    16'd1375: out <= 16'hFDBE;
    16'd1376: out <= 16'h03C6;    16'd1377: out <= 16'h0132;    16'd1378: out <= 16'h0400;    16'd1379: out <= 16'h0434;
    16'd1380: out <= 16'h06F0;    16'd1381: out <= 16'hFD77;    16'd1382: out <= 16'hFD50;    16'd1383: out <= 16'hFD84;
    16'd1384: out <= 16'hFD44;    16'd1385: out <= 16'hFDB5;    16'd1386: out <= 16'h054B;    16'd1387: out <= 16'hFF21;
    16'd1388: out <= 16'h0026;    16'd1389: out <= 16'h0164;    16'd1390: out <= 16'hFD0A;    16'd1391: out <= 16'h0019;
    16'd1392: out <= 16'h04D7;    16'd1393: out <= 16'h01C2;    16'd1394: out <= 16'h0200;    16'd1395: out <= 16'h06AA;
    16'd1396: out <= 16'hFF49;    16'd1397: out <= 16'h02FF;    16'd1398: out <= 16'hFEC3;    16'd1399: out <= 16'hFDC0;
    16'd1400: out <= 16'h031E;    16'd1401: out <= 16'h0844;    16'd1402: out <= 16'h0421;    16'd1403: out <= 16'h060E;
    16'd1404: out <= 16'h0525;    16'd1405: out <= 16'hF9CB;    16'd1406: out <= 16'h0516;    16'd1407: out <= 16'h062D;
    16'd1408: out <= 16'hFFC4;    16'd1409: out <= 16'hFFF0;    16'd1410: out <= 16'hFBDC;    16'd1411: out <= 16'hFFFB;
    16'd1412: out <= 16'h01A9;    16'd1413: out <= 16'hFD39;    16'd1414: out <= 16'hF813;    16'd1415: out <= 16'h0251;
    16'd1416: out <= 16'h0726;    16'd1417: out <= 16'h00C1;    16'd1418: out <= 16'hFF85;    16'd1419: out <= 16'hFA06;
    16'd1420: out <= 16'hF707;    16'd1421: out <= 16'h01DB;    16'd1422: out <= 16'hFF54;    16'd1423: out <= 16'h00D4;
    16'd1424: out <= 16'h0189;    16'd1425: out <= 16'hFF4E;    16'd1426: out <= 16'h05C2;    16'd1427: out <= 16'h03C0;
    16'd1428: out <= 16'h05F9;    16'd1429: out <= 16'hFF9F;    16'd1430: out <= 16'hFEB6;    16'd1431: out <= 16'h0033;
    16'd1432: out <= 16'hFC8D;    16'd1433: out <= 16'h015F;    16'd1434: out <= 16'hFD8C;    16'd1435: out <= 16'hFC71;
    16'd1436: out <= 16'h0246;    16'd1437: out <= 16'hFAEB;    16'd1438: out <= 16'h0978;    16'd1439: out <= 16'hF5EE;
    16'd1440: out <= 16'h082C;    16'd1441: out <= 16'hFE64;    16'd1442: out <= 16'h005E;    16'd1443: out <= 16'hFE11;
    16'd1444: out <= 16'hFE2E;    16'd1445: out <= 16'h028B;    16'd1446: out <= 16'h02D5;    16'd1447: out <= 16'h053B;
    16'd1448: out <= 16'hFA3B;    16'd1449: out <= 16'hFEEC;    16'd1450: out <= 16'hFBD9;    16'd1451: out <= 16'hF9BF;
    16'd1452: out <= 16'hFD00;    16'd1453: out <= 16'hFFF9;    16'd1454: out <= 16'hFDF7;    16'd1455: out <= 16'h0728;
    16'd1456: out <= 16'hFC40;    16'd1457: out <= 16'hFE95;    16'd1458: out <= 16'h00BD;    16'd1459: out <= 16'hFF83;
    16'd1460: out <= 16'hFB78;    16'd1461: out <= 16'h030B;    16'd1462: out <= 16'h0508;    16'd1463: out <= 16'hF878;
    16'd1464: out <= 16'hFEAD;    16'd1465: out <= 16'hFEA3;    16'd1466: out <= 16'h00A6;    16'd1467: out <= 16'hFF50;
    16'd1468: out <= 16'h05B1;    16'd1469: out <= 16'hFF95;    16'd1470: out <= 16'h03A9;    16'd1471: out <= 16'h01C1;
    16'd1472: out <= 16'hFE13;    16'd1473: out <= 16'h01C3;    16'd1474: out <= 16'h00B3;    16'd1475: out <= 16'h04A4;
    16'd1476: out <= 16'hFC0C;    16'd1477: out <= 16'h0264;    16'd1478: out <= 16'hFB0F;    16'd1479: out <= 16'h0013;
    16'd1480: out <= 16'h049F;    16'd1481: out <= 16'hF9FD;    16'd1482: out <= 16'hFCDA;    16'd1483: out <= 16'hFEDD;
    16'd1484: out <= 16'h05C0;    16'd1485: out <= 16'h05B5;    16'd1486: out <= 16'h06D8;    16'd1487: out <= 16'hFED0;
    16'd1488: out <= 16'hFF4D;    16'd1489: out <= 16'h0239;    16'd1490: out <= 16'hFAD5;    16'd1491: out <= 16'h031D;
    16'd1492: out <= 16'h043E;    16'd1493: out <= 16'hFA0E;    16'd1494: out <= 16'h0096;    16'd1495: out <= 16'h0178;
    16'd1496: out <= 16'hFFAD;    16'd1497: out <= 16'hFF5E;    16'd1498: out <= 16'hFBC2;    16'd1499: out <= 16'h03E9;
    16'd1500: out <= 16'hFC9E;    16'd1501: out <= 16'h0091;    16'd1502: out <= 16'h0591;    16'd1503: out <= 16'hFEC6;
    16'd1504: out <= 16'hFBF6;    16'd1505: out <= 16'hFE84;    16'd1506: out <= 16'h008A;    16'd1507: out <= 16'h04CB;
    16'd1508: out <= 16'hFC7C;    16'd1509: out <= 16'h04EC;    16'd1510: out <= 16'h0084;    16'd1511: out <= 16'h0348;
    16'd1512: out <= 16'h03DF;    16'd1513: out <= 16'h002F;    16'd1514: out <= 16'h04C0;    16'd1515: out <= 16'h00FF;
    16'd1516: out <= 16'hFE4A;    16'd1517: out <= 16'h03DF;    16'd1518: out <= 16'hFD61;    16'd1519: out <= 16'h06D2;
    16'd1520: out <= 16'hFB7F;    16'd1521: out <= 16'hF8B5;    16'd1522: out <= 16'hFDD6;    16'd1523: out <= 16'hFF47;
    16'd1524: out <= 16'h03B4;    16'd1525: out <= 16'hFA7C;    16'd1526: out <= 16'hFC56;    16'd1527: out <= 16'hF94E;
    16'd1528: out <= 16'hF54E;    16'd1529: out <= 16'hFA4E;    16'd1530: out <= 16'hFA7A;    16'd1531: out <= 16'h0538;
    16'd1532: out <= 16'h0323;    16'd1533: out <= 16'hFAE8;    16'd1534: out <= 16'h0010;    16'd1535: out <= 16'h00A9;
    16'd1536: out <= 16'hFF21;    16'd1537: out <= 16'hFC12;    16'd1538: out <= 16'hFBF5;    16'd1539: out <= 16'h00BF;
    16'd1540: out <= 16'h00EA;    16'd1541: out <= 16'hFDC9;    16'd1542: out <= 16'h00F1;    16'd1543: out <= 16'h06E5;
    16'd1544: out <= 16'hFFD2;    16'd1545: out <= 16'hF8A7;    16'd1546: out <= 16'h0118;    16'd1547: out <= 16'h08EB;
    16'd1548: out <= 16'hF944;    16'd1549: out <= 16'hFA2C;    16'd1550: out <= 16'h00A8;    16'd1551: out <= 16'hFFA8;
    16'd1552: out <= 16'hFFFB;    16'd1553: out <= 16'hFE8A;    16'd1554: out <= 16'h0202;    16'd1555: out <= 16'hFAD6;
    16'd1556: out <= 16'hFA04;    16'd1557: out <= 16'h0254;    16'd1558: out <= 16'h0827;    16'd1559: out <= 16'h008F;
    16'd1560: out <= 16'hFB15;    16'd1561: out <= 16'hFAF1;    16'd1562: out <= 16'h005F;    16'd1563: out <= 16'h0306;
    16'd1564: out <= 16'h02D4;    16'd1565: out <= 16'hFB6D;    16'd1566: out <= 16'h00F3;    16'd1567: out <= 16'h04CC;
    16'd1568: out <= 16'h069B;    16'd1569: out <= 16'h006F;    16'd1570: out <= 16'hFBBB;    16'd1571: out <= 16'h08DD;
    16'd1572: out <= 16'h0290;    16'd1573: out <= 16'hFC29;    16'd1574: out <= 16'h0399;    16'd1575: out <= 16'h01C2;
    16'd1576: out <= 16'h0167;    16'd1577: out <= 16'h0D0C;    16'd1578: out <= 16'hFE3F;    16'd1579: out <= 16'hFFF4;
    16'd1580: out <= 16'hFD1C;    16'd1581: out <= 16'h0118;    16'd1582: out <= 16'h001A;    16'd1583: out <= 16'hFCAC;
    16'd1584: out <= 16'hFE89;    16'd1585: out <= 16'h011A;    16'd1586: out <= 16'hFAB0;    16'd1587: out <= 16'hFF49;
    16'd1588: out <= 16'h03B5;    16'd1589: out <= 16'hFC67;    16'd1590: out <= 16'hFED9;    16'd1591: out <= 16'h0141;
    16'd1592: out <= 16'h0204;    16'd1593: out <= 16'hFFE6;    16'd1594: out <= 16'h005D;    16'd1595: out <= 16'hFD89;
    16'd1596: out <= 16'h0059;    16'd1597: out <= 16'hFF7F;    16'd1598: out <= 16'hFC33;    16'd1599: out <= 16'hFC1B;
    16'd1600: out <= 16'hFB0A;    16'd1601: out <= 16'hFCD3;    16'd1602: out <= 16'h01DF;    16'd1603: out <= 16'h0306;
    16'd1604: out <= 16'hF7AE;    16'd1605: out <= 16'hFCAC;    16'd1606: out <= 16'h06D0;    16'd1607: out <= 16'h02C6;
    16'd1608: out <= 16'h0722;    16'd1609: out <= 16'h08D7;    16'd1610: out <= 16'h0436;    16'd1611: out <= 16'hF8CF;
    16'd1612: out <= 16'hFFA7;    16'd1613: out <= 16'h020E;    16'd1614: out <= 16'h0277;    16'd1615: out <= 16'hFD40;
    16'd1616: out <= 16'h0312;    16'd1617: out <= 16'hFE7F;    16'd1618: out <= 16'hFD34;    16'd1619: out <= 16'h01CE;
    16'd1620: out <= 16'h05D0;    16'd1621: out <= 16'hFD85;    16'd1622: out <= 16'h0094;    16'd1623: out <= 16'hFA0F;
    16'd1624: out <= 16'hFFC5;    16'd1625: out <= 16'h0661;    16'd1626: out <= 16'h08A7;    16'd1627: out <= 16'hFE75;
    16'd1628: out <= 16'h009E;    16'd1629: out <= 16'hFEC7;    16'd1630: out <= 16'h0387;    16'd1631: out <= 16'h0249;
    16'd1632: out <= 16'h030E;    16'd1633: out <= 16'h0439;    16'd1634: out <= 16'hFFC6;    16'd1635: out <= 16'hFCF5;
    16'd1636: out <= 16'hFCAB;    16'd1637: out <= 16'hFF42;    16'd1638: out <= 16'h040E;    16'd1639: out <= 16'hFBFD;
    16'd1640: out <= 16'h0334;    16'd1641: out <= 16'hFB6E;    16'd1642: out <= 16'hFE16;    16'd1643: out <= 16'h0191;
    16'd1644: out <= 16'h01A5;    16'd1645: out <= 16'hFF2B;    16'd1646: out <= 16'h0559;    16'd1647: out <= 16'hFF81;
    16'd1648: out <= 16'hF798;    16'd1649: out <= 16'h0062;    16'd1650: out <= 16'h01B2;    16'd1651: out <= 16'h0A0B;
    16'd1652: out <= 16'hFE05;    16'd1653: out <= 16'h005E;    16'd1654: out <= 16'h038F;    16'd1655: out <= 16'h0243;
    16'd1656: out <= 16'h06AB;    16'd1657: out <= 16'hF972;    16'd1658: out <= 16'h006E;    16'd1659: out <= 16'h01E5;
    16'd1660: out <= 16'h05E1;    16'd1661: out <= 16'hFDC7;    16'd1662: out <= 16'h0648;    16'd1663: out <= 16'hFCD4;
    16'd1664: out <= 16'hFD7B;    16'd1665: out <= 16'h001E;    16'd1666: out <= 16'h04D7;    16'd1667: out <= 16'hFD8E;
    16'd1668: out <= 16'hFB5C;    16'd1669: out <= 16'hFA21;    16'd1670: out <= 16'hFCBB;    16'd1671: out <= 16'hFC24;
    16'd1672: out <= 16'h0347;    16'd1673: out <= 16'h01E4;    16'd1674: out <= 16'hFBD5;    16'd1675: out <= 16'hF92F;
    16'd1676: out <= 16'h0052;    16'd1677: out <= 16'h07E2;    16'd1678: out <= 16'hFBCB;    16'd1679: out <= 16'h093A;
    16'd1680: out <= 16'h021C;    16'd1681: out <= 16'h031C;    16'd1682: out <= 16'hFB85;    16'd1683: out <= 16'hF50F;
    16'd1684: out <= 16'h061A;    16'd1685: out <= 16'hFAD0;    16'd1686: out <= 16'hF60F;    16'd1687: out <= 16'hFF25;
    16'd1688: out <= 16'h028C;    16'd1689: out <= 16'hFCCF;    16'd1690: out <= 16'hFE00;    16'd1691: out <= 16'h05D7;
    16'd1692: out <= 16'hFA8E;    16'd1693: out <= 16'h03BC;    16'd1694: out <= 16'h02AF;    16'd1695: out <= 16'h00F4;
    16'd1696: out <= 16'h05DA;    16'd1697: out <= 16'h050F;    16'd1698: out <= 16'h00FB;    16'd1699: out <= 16'hFFD5;
    16'd1700: out <= 16'hFFBB;    16'd1701: out <= 16'hFE0F;    16'd1702: out <= 16'hFE6E;    16'd1703: out <= 16'hFF8A;
    16'd1704: out <= 16'h04E7;    16'd1705: out <= 16'hFB32;    16'd1706: out <= 16'h01A4;    16'd1707: out <= 16'hFFD0;
    16'd1708: out <= 16'hFE12;    16'd1709: out <= 16'h0290;    16'd1710: out <= 16'h01C4;    16'd1711: out <= 16'h01EC;
    16'd1712: out <= 16'hFD83;    16'd1713: out <= 16'hFD98;    16'd1714: out <= 16'h01CB;    16'd1715: out <= 16'hFB26;
    16'd1716: out <= 16'hFF9E;    16'd1717: out <= 16'hFBCE;    16'd1718: out <= 16'hFE46;    16'd1719: out <= 16'hFAC4;
    16'd1720: out <= 16'hFE37;    16'd1721: out <= 16'hFEB2;    16'd1722: out <= 16'hFB7F;    16'd1723: out <= 16'h01B3;
    16'd1724: out <= 16'hFFDF;    16'd1725: out <= 16'h0424;    16'd1726: out <= 16'hFB6B;    16'd1727: out <= 16'h0448;
    16'd1728: out <= 16'hFA8B;    16'd1729: out <= 16'hFC58;    16'd1730: out <= 16'hFD5B;    16'd1731: out <= 16'hFECA;
    16'd1732: out <= 16'hFC02;    16'd1733: out <= 16'h0271;    16'd1734: out <= 16'hF9F1;    16'd1735: out <= 16'hFA30;
    16'd1736: out <= 16'hFFE4;    16'd1737: out <= 16'h04BB;    16'd1738: out <= 16'h008E;    16'd1739: out <= 16'h01A4;
    16'd1740: out <= 16'h021C;    16'd1741: out <= 16'hFDF1;    16'd1742: out <= 16'h00E7;    16'd1743: out <= 16'h008F;
    16'd1744: out <= 16'hF8FA;    16'd1745: out <= 16'hF953;    16'd1746: out <= 16'h032F;    16'd1747: out <= 16'hFC0A;
    16'd1748: out <= 16'hF980;    16'd1749: out <= 16'hFE52;    16'd1750: out <= 16'h0309;    16'd1751: out <= 16'h01B3;
    16'd1752: out <= 16'h05D0;    16'd1753: out <= 16'h0388;    16'd1754: out <= 16'hFE51;    16'd1755: out <= 16'h0247;
    16'd1756: out <= 16'hFAF1;    16'd1757: out <= 16'hFE78;    16'd1758: out <= 16'hFFD5;    16'd1759: out <= 16'h001E;
    16'd1760: out <= 16'h0505;    16'd1761: out <= 16'h04CF;    16'd1762: out <= 16'h0070;    16'd1763: out <= 16'hFC89;
    16'd1764: out <= 16'h0326;    16'd1765: out <= 16'hFE66;    16'd1766: out <= 16'h00AA;    16'd1767: out <= 16'h0041;
    16'd1768: out <= 16'h035D;    16'd1769: out <= 16'h028C;    16'd1770: out <= 16'hFE09;    16'd1771: out <= 16'h04CD;
    16'd1772: out <= 16'h031C;    16'd1773: out <= 16'h00A9;    16'd1774: out <= 16'hFFCF;    16'd1775: out <= 16'h0470;
    16'd1776: out <= 16'h007F;    16'd1777: out <= 16'h01F5;    16'd1778: out <= 16'h030E;    16'd1779: out <= 16'hFF42;
    16'd1780: out <= 16'h01E2;    16'd1781: out <= 16'hFAD8;    16'd1782: out <= 16'h0103;    16'd1783: out <= 16'hFE67;
    16'd1784: out <= 16'hFE93;    16'd1785: out <= 16'hFD74;    16'd1786: out <= 16'h0056;    16'd1787: out <= 16'hFFF8;
    16'd1788: out <= 16'h02A0;    16'd1789: out <= 16'hFB77;    16'd1790: out <= 16'h03E1;    16'd1791: out <= 16'hFEAC;
    16'd1792: out <= 16'h0533;    16'd1793: out <= 16'hFE32;    16'd1794: out <= 16'h0247;    16'd1795: out <= 16'hFF0F;
    16'd1796: out <= 16'h0075;    16'd1797: out <= 16'h01E3;    16'd1798: out <= 16'hFC9C;    16'd1799: out <= 16'hFB5B;
    16'd1800: out <= 16'hF836;    16'd1801: out <= 16'h043C;    16'd1802: out <= 16'h020A;    16'd1803: out <= 16'h04DE;
    16'd1804: out <= 16'hFBF7;    16'd1805: out <= 16'hFC77;    16'd1806: out <= 16'hF9BB;    16'd1807: out <= 16'h01DC;
    16'd1808: out <= 16'hFC56;    16'd1809: out <= 16'hFD7D;    16'd1810: out <= 16'hFE25;    16'd1811: out <= 16'hF9B3;
    16'd1812: out <= 16'h0777;    16'd1813: out <= 16'h046F;    16'd1814: out <= 16'hFD4A;    16'd1815: out <= 16'h026F;
    16'd1816: out <= 16'h0259;    16'd1817: out <= 16'hFA37;    16'd1818: out <= 16'hFD9C;    16'd1819: out <= 16'hFF26;
    16'd1820: out <= 16'hFF8D;    16'd1821: out <= 16'h0149;    16'd1822: out <= 16'hFAEE;    16'd1823: out <= 16'hFDB8;
    16'd1824: out <= 16'h0274;    16'd1825: out <= 16'h0267;    16'd1826: out <= 16'h013A;    16'd1827: out <= 16'h0626;
    16'd1828: out <= 16'hFB23;    16'd1829: out <= 16'h010A;    16'd1830: out <= 16'h0890;    16'd1831: out <= 16'hFC0F;
    16'd1832: out <= 16'hFCF3;    16'd1833: out <= 16'h04E4;    16'd1834: out <= 16'hF8E0;    16'd1835: out <= 16'hFB1C;
    16'd1836: out <= 16'hFFE6;    16'd1837: out <= 16'h0A41;    16'd1838: out <= 16'h06FE;    16'd1839: out <= 16'hFEB3;
    16'd1840: out <= 16'hFBF1;    16'd1841: out <= 16'h0541;    16'd1842: out <= 16'hFDF5;    16'd1843: out <= 16'h0493;
    16'd1844: out <= 16'hF7D2;    16'd1845: out <= 16'h0907;    16'd1846: out <= 16'h0152;    16'd1847: out <= 16'hFD4E;
    16'd1848: out <= 16'h084E;    16'd1849: out <= 16'h061B;    16'd1850: out <= 16'hFAE4;    16'd1851: out <= 16'h0421;
    16'd1852: out <= 16'hF827;    16'd1853: out <= 16'hFBAC;    16'd1854: out <= 16'h02DE;    16'd1855: out <= 16'h0418;
    16'd1856: out <= 16'hFE04;    16'd1857: out <= 16'hFE5C;    16'd1858: out <= 16'h0894;    16'd1859: out <= 16'h0162;
    16'd1860: out <= 16'h0043;    16'd1861: out <= 16'hFD04;    16'd1862: out <= 16'hFA0E;    16'd1863: out <= 16'h00E8;
    16'd1864: out <= 16'h011B;    16'd1865: out <= 16'h0440;    16'd1866: out <= 16'h0292;    16'd1867: out <= 16'hF95E;
    16'd1868: out <= 16'h0A28;    16'd1869: out <= 16'h08BD;    16'd1870: out <= 16'h039E;    16'd1871: out <= 16'h0094;
    16'd1872: out <= 16'h007E;    16'd1873: out <= 16'hFD31;    16'd1874: out <= 16'hFB9F;    16'd1875: out <= 16'hFD33;
    16'd1876: out <= 16'h0063;    16'd1877: out <= 16'h0383;    16'd1878: out <= 16'hFCEC;    16'd1879: out <= 16'hFACD;
    16'd1880: out <= 16'h0A2E;    16'd1881: out <= 16'hFC4A;    16'd1882: out <= 16'h0148;    16'd1883: out <= 16'h0381;
    16'd1884: out <= 16'h01B6;    16'd1885: out <= 16'h0195;    16'd1886: out <= 16'h0153;    16'd1887: out <= 16'hFD41;
    16'd1888: out <= 16'h0713;    16'd1889: out <= 16'h06DD;    16'd1890: out <= 16'h0413;    16'd1891: out <= 16'hFCCB;
    16'd1892: out <= 16'hFEC0;    16'd1893: out <= 16'hFE30;    16'd1894: out <= 16'h0334;    16'd1895: out <= 16'hFF54;
    16'd1896: out <= 16'h0353;    16'd1897: out <= 16'hFE2C;    16'd1898: out <= 16'hFC0E;    16'd1899: out <= 16'hFBF4;
    16'd1900: out <= 16'h0035;    16'd1901: out <= 16'h059A;    16'd1902: out <= 16'h0402;    16'd1903: out <= 16'hFAD4;
    16'd1904: out <= 16'h009D;    16'd1905: out <= 16'hFC4F;    16'd1906: out <= 16'hFE9B;    16'd1907: out <= 16'hFF37;
    16'd1908: out <= 16'hF9A9;    16'd1909: out <= 16'h01FA;    16'd1910: out <= 16'hFDC7;    16'd1911: out <= 16'hFD42;
    16'd1912: out <= 16'hFE06;    16'd1913: out <= 16'h03DA;    16'd1914: out <= 16'h082C;    16'd1915: out <= 16'h005E;
    16'd1916: out <= 16'hFC47;    16'd1917: out <= 16'h0476;    16'd1918: out <= 16'hFA2D;    16'd1919: out <= 16'hFD05;
    16'd1920: out <= 16'h0618;    16'd1921: out <= 16'h0320;    16'd1922: out <= 16'hFF1B;    16'd1923: out <= 16'h05B5;
    16'd1924: out <= 16'h008A;    16'd1925: out <= 16'h0029;    16'd1926: out <= 16'hFD6D;    16'd1927: out <= 16'hFF05;
    16'd1928: out <= 16'hFF85;    16'd1929: out <= 16'hFE0A;    16'd1930: out <= 16'hFF59;    16'd1931: out <= 16'h025A;
    16'd1932: out <= 16'h0012;    16'd1933: out <= 16'h00BB;    16'd1934: out <= 16'hFAAE;    16'd1935: out <= 16'hFC90;
    16'd1936: out <= 16'h06E2;    16'd1937: out <= 16'hFDA4;    16'd1938: out <= 16'hFDE5;    16'd1939: out <= 16'h07B7;
    16'd1940: out <= 16'hFA32;    16'd1941: out <= 16'h062F;    16'd1942: out <= 16'hFABE;    16'd1943: out <= 16'hFDEE;
    16'd1944: out <= 16'h0169;    16'd1945: out <= 16'hFEC5;    16'd1946: out <= 16'hFA3E;    16'd1947: out <= 16'hFF26;
    16'd1948: out <= 16'h00D4;    16'd1949: out <= 16'hFE61;    16'd1950: out <= 16'hFD15;    16'd1951: out <= 16'hFDDF;
    16'd1952: out <= 16'hFF8F;    16'd1953: out <= 16'h00ED;    16'd1954: out <= 16'h00AA;    16'd1955: out <= 16'hFE7E;
    16'd1956: out <= 16'h030A;    16'd1957: out <= 16'h094D;    16'd1958: out <= 16'hFC95;    16'd1959: out <= 16'hFFBA;
    16'd1960: out <= 16'h023A;    16'd1961: out <= 16'h043D;    16'd1962: out <= 16'h0469;    16'd1963: out <= 16'h00A7;
    16'd1964: out <= 16'h037F;    16'd1965: out <= 16'hFC47;    16'd1966: out <= 16'h0024;    16'd1967: out <= 16'hFA07;
    16'd1968: out <= 16'hFF1F;    16'd1969: out <= 16'h02AD;    16'd1970: out <= 16'h01EF;    16'd1971: out <= 16'h0452;
    16'd1972: out <= 16'h05F1;    16'd1973: out <= 16'h03E6;    16'd1974: out <= 16'hFDB2;    16'd1975: out <= 16'h003D;
    16'd1976: out <= 16'hFB23;    16'd1977: out <= 16'h079F;    16'd1978: out <= 16'h0156;    16'd1979: out <= 16'hFF44;
    16'd1980: out <= 16'h0399;    16'd1981: out <= 16'hFE3C;    16'd1982: out <= 16'h014A;    16'd1983: out <= 16'hFAF7;
    16'd1984: out <= 16'hFFDD;    16'd1985: out <= 16'h030F;    16'd1986: out <= 16'hFF58;    16'd1987: out <= 16'h008A;
    16'd1988: out <= 16'hFDF8;    16'd1989: out <= 16'h02E0;    16'd1990: out <= 16'h0484;    16'd1991: out <= 16'h01FB;
    16'd1992: out <= 16'hFEE4;    16'd1993: out <= 16'hFD1B;    16'd1994: out <= 16'hF98F;    16'd1995: out <= 16'h0112;
    16'd1996: out <= 16'hFC9E;    16'd1997: out <= 16'h04FB;    16'd1998: out <= 16'hFE6B;    16'd1999: out <= 16'hFF6F;
    16'd2000: out <= 16'hF914;    16'd2001: out <= 16'hFB21;    16'd2002: out <= 16'hFCE1;    16'd2003: out <= 16'hF968;
    16'd2004: out <= 16'h0126;    16'd2005: out <= 16'hFBC5;    16'd2006: out <= 16'hFC1F;    16'd2007: out <= 16'hF8BE;
    16'd2008: out <= 16'h04B1;    16'd2009: out <= 16'h05AF;    16'd2010: out <= 16'hFCF8;    16'd2011: out <= 16'h0257;
    16'd2012: out <= 16'hFEF9;    16'd2013: out <= 16'hFFEB;    16'd2014: out <= 16'hFB84;    16'd2015: out <= 16'h003B;
    16'd2016: out <= 16'h04C0;    16'd2017: out <= 16'hF826;    16'd2018: out <= 16'h0019;    16'd2019: out <= 16'hFB23;
    16'd2020: out <= 16'hFEF7;    16'd2021: out <= 16'h007E;    16'd2022: out <= 16'h0054;    16'd2023: out <= 16'h0343;
    16'd2024: out <= 16'h057B;    16'd2025: out <= 16'hFCCA;    16'd2026: out <= 16'h028F;    16'd2027: out <= 16'h097F;
    16'd2028: out <= 16'h015A;    16'd2029: out <= 16'h02F7;    16'd2030: out <= 16'h0372;    16'd2031: out <= 16'h0698;
    16'd2032: out <= 16'h021A;    16'd2033: out <= 16'h02C7;    16'd2034: out <= 16'hFC87;    16'd2035: out <= 16'h0346;
    16'd2036: out <= 16'hF822;    16'd2037: out <= 16'hFB5D;    16'd2038: out <= 16'h05C9;    16'd2039: out <= 16'h0009;
    16'd2040: out <= 16'h0324;    16'd2041: out <= 16'hFF81;    16'd2042: out <= 16'hFFB3;    16'd2043: out <= 16'h014B;
    16'd2044: out <= 16'hFEA0;    16'd2045: out <= 16'h03A8;    16'd2046: out <= 16'hFE2B;    16'd2047: out <= 16'h00A5;
    16'd2048: out <= 16'h00A9;    16'd2049: out <= 16'h026D;    16'd2050: out <= 16'hFE6F;    16'd2051: out <= 16'h006D;
    16'd2052: out <= 16'h0944;    16'd2053: out <= 16'hFB8E;    16'd2054: out <= 16'hFD11;    16'd2055: out <= 16'h040A;
    16'd2056: out <= 16'hFB66;    16'd2057: out <= 16'h026B;    16'd2058: out <= 16'h0008;    16'd2059: out <= 16'h046F;
    16'd2060: out <= 16'hF8AD;    16'd2061: out <= 16'hFC28;    16'd2062: out <= 16'hFF04;    16'd2063: out <= 16'hFEF8;
    16'd2064: out <= 16'h04FF;    16'd2065: out <= 16'h0670;    16'd2066: out <= 16'hF68A;    16'd2067: out <= 16'h0587;
    16'd2068: out <= 16'h00E1;    16'd2069: out <= 16'hFCF0;    16'd2070: out <= 16'h0051;    16'd2071: out <= 16'hFB91;
    16'd2072: out <= 16'h03C9;    16'd2073: out <= 16'h0464;    16'd2074: out <= 16'h0780;    16'd2075: out <= 16'h03C4;
    16'd2076: out <= 16'h0015;    16'd2077: out <= 16'hF858;    16'd2078: out <= 16'h0830;    16'd2079: out <= 16'hFB45;
    16'd2080: out <= 16'hFE96;    16'd2081: out <= 16'h0308;    16'd2082: out <= 16'hFF4B;    16'd2083: out <= 16'hFD58;
    16'd2084: out <= 16'hFC28;    16'd2085: out <= 16'h0196;    16'd2086: out <= 16'h0622;    16'd2087: out <= 16'hFFB6;
    16'd2088: out <= 16'h003F;    16'd2089: out <= 16'h030A;    16'd2090: out <= 16'hFDBA;    16'd2091: out <= 16'hFAB1;
    16'd2092: out <= 16'hFF03;    16'd2093: out <= 16'h021C;    16'd2094: out <= 16'hFE84;    16'd2095: out <= 16'hFE9A;
    16'd2096: out <= 16'h0086;    16'd2097: out <= 16'hFFAC;    16'd2098: out <= 16'h009F;    16'd2099: out <= 16'hFE81;
    16'd2100: out <= 16'h005E;    16'd2101: out <= 16'h0440;    16'd2102: out <= 16'h0194;    16'd2103: out <= 16'hFF83;
    16'd2104: out <= 16'hFE0F;    16'd2105: out <= 16'h0191;    16'd2106: out <= 16'hFCF4;    16'd2107: out <= 16'hFB61;
    16'd2108: out <= 16'h038A;    16'd2109: out <= 16'hF8E9;    16'd2110: out <= 16'h021E;    16'd2111: out <= 16'hFDCE;
    16'd2112: out <= 16'h028A;    16'd2113: out <= 16'h0633;    16'd2114: out <= 16'h07EB;    16'd2115: out <= 16'h0B3A;
    16'd2116: out <= 16'hFFBC;    16'd2117: out <= 16'h02A1;    16'd2118: out <= 16'h0808;    16'd2119: out <= 16'hFE95;
    16'd2120: out <= 16'h03A3;    16'd2121: out <= 16'h036B;    16'd2122: out <= 16'hFCD9;    16'd2123: out <= 16'h019C;
    16'd2124: out <= 16'h0776;    16'd2125: out <= 16'h0139;    16'd2126: out <= 16'h03B7;    16'd2127: out <= 16'hFEA0;
    16'd2128: out <= 16'h05A7;    16'd2129: out <= 16'hFDC7;    16'd2130: out <= 16'hF9FE;    16'd2131: out <= 16'h034F;
    16'd2132: out <= 16'hFC20;    16'd2133: out <= 16'hFAFD;    16'd2134: out <= 16'h004D;    16'd2135: out <= 16'hFCD8;
    16'd2136: out <= 16'hFFAA;    16'd2137: out <= 16'hFC9E;    16'd2138: out <= 16'h0665;    16'd2139: out <= 16'hFB4B;
    16'd2140: out <= 16'h0011;    16'd2141: out <= 16'hFA4B;    16'd2142: out <= 16'hFCA9;    16'd2143: out <= 16'h024C;
    16'd2144: out <= 16'hFEF7;    16'd2145: out <= 16'hFF1B;    16'd2146: out <= 16'hFE62;    16'd2147: out <= 16'hFF2A;
    16'd2148: out <= 16'h0213;    16'd2149: out <= 16'hFC1C;    16'd2150: out <= 16'hFD7F;    16'd2151: out <= 16'hFE8F;
    16'd2152: out <= 16'hFE11;    16'd2153: out <= 16'hFFB4;    16'd2154: out <= 16'hFD30;    16'd2155: out <= 16'h01AB;
    16'd2156: out <= 16'h01A2;    16'd2157: out <= 16'hFB98;    16'd2158: out <= 16'hFAB3;    16'd2159: out <= 16'hFCCE;
    16'd2160: out <= 16'hFA7B;    16'd2161: out <= 16'h052A;    16'd2162: out <= 16'h00C7;    16'd2163: out <= 16'hFF9F;
    16'd2164: out <= 16'h00F5;    16'd2165: out <= 16'h006F;    16'd2166: out <= 16'h00B3;    16'd2167: out <= 16'hFBC0;
    16'd2168: out <= 16'hFC52;    16'd2169: out <= 16'h04BF;    16'd2170: out <= 16'hFF5E;    16'd2171: out <= 16'hFDED;
    16'd2172: out <= 16'h04D0;    16'd2173: out <= 16'hFCB7;    16'd2174: out <= 16'hFEB0;    16'd2175: out <= 16'h03C3;
    16'd2176: out <= 16'h04D3;    16'd2177: out <= 16'h0291;    16'd2178: out <= 16'h00B8;    16'd2179: out <= 16'h034B;
    16'd2180: out <= 16'hFD48;    16'd2181: out <= 16'h0197;    16'd2182: out <= 16'h0612;    16'd2183: out <= 16'hFD9A;
    16'd2184: out <= 16'hFDC2;    16'd2185: out <= 16'hFA58;    16'd2186: out <= 16'hFF06;    16'd2187: out <= 16'h03EC;
    16'd2188: out <= 16'h00F8;    16'd2189: out <= 16'h050E;    16'd2190: out <= 16'h00D1;    16'd2191: out <= 16'hFD7D;
    16'd2192: out <= 16'h054A;    16'd2193: out <= 16'hFF8D;    16'd2194: out <= 16'h00D9;    16'd2195: out <= 16'hFFE5;
    16'd2196: out <= 16'h07B3;    16'd2197: out <= 16'h05F5;    16'd2198: out <= 16'hFC49;    16'd2199: out <= 16'h0344;
    16'd2200: out <= 16'h0479;    16'd2201: out <= 16'h03B1;    16'd2202: out <= 16'h01CC;    16'd2203: out <= 16'h000F;
    16'd2204: out <= 16'h0116;    16'd2205: out <= 16'hFFDB;    16'd2206: out <= 16'hFFF1;    16'd2207: out <= 16'hF8F2;
    16'd2208: out <= 16'hFB37;    16'd2209: out <= 16'hFCB3;    16'd2210: out <= 16'hFEB0;    16'd2211: out <= 16'h05A1;
    16'd2212: out <= 16'hFD79;    16'd2213: out <= 16'h0192;    16'd2214: out <= 16'hFECC;    16'd2215: out <= 16'h0013;
    16'd2216: out <= 16'hFACB;    16'd2217: out <= 16'hFFA5;    16'd2218: out <= 16'hFFA0;    16'd2219: out <= 16'h00F4;
    16'd2220: out <= 16'h0306;    16'd2221: out <= 16'hFE20;    16'd2222: out <= 16'hFE8E;    16'd2223: out <= 16'hFD61;
    16'd2224: out <= 16'hFBD8;    16'd2225: out <= 16'hFED9;    16'd2226: out <= 16'h02BD;    16'd2227: out <= 16'h00CF;
    16'd2228: out <= 16'hF949;    16'd2229: out <= 16'hFBCD;    16'd2230: out <= 16'hFF43;    16'd2231: out <= 16'hFE0B;
    16'd2232: out <= 16'h01FD;    16'd2233: out <= 16'hFA36;    16'd2234: out <= 16'hFB68;    16'd2235: out <= 16'h00E2;
    16'd2236: out <= 16'hFF8F;    16'd2237: out <= 16'h0148;    16'd2238: out <= 16'h0059;    16'd2239: out <= 16'hF906;
    16'd2240: out <= 16'h0168;    16'd2241: out <= 16'h02D3;    16'd2242: out <= 16'hFEA9;    16'd2243: out <= 16'hFE64;
    16'd2244: out <= 16'hFCC3;    16'd2245: out <= 16'hFAE9;    16'd2246: out <= 16'h04BB;    16'd2247: out <= 16'h0143;
    16'd2248: out <= 16'hFE66;    16'd2249: out <= 16'hFF76;    16'd2250: out <= 16'hFFFB;    16'd2251: out <= 16'h0294;
    16'd2252: out <= 16'hFF4B;    16'd2253: out <= 16'h044F;    16'd2254: out <= 16'hFADB;    16'd2255: out <= 16'h0284;
    16'd2256: out <= 16'h069A;    16'd2257: out <= 16'hFD88;    16'd2258: out <= 16'hFBD7;    16'd2259: out <= 16'hFEB4;
    16'd2260: out <= 16'hFFAB;    16'd2261: out <= 16'hFB5D;    16'd2262: out <= 16'hFF69;    16'd2263: out <= 16'h013D;
    16'd2264: out <= 16'hFD47;    16'd2265: out <= 16'hFAD7;    16'd2266: out <= 16'h026F;    16'd2267: out <= 16'hFF68;
    16'd2268: out <= 16'hFDE5;    16'd2269: out <= 16'h027C;    16'd2270: out <= 16'hFF23;    16'd2271: out <= 16'hF639;
    16'd2272: out <= 16'hFAA5;    16'd2273: out <= 16'h0354;    16'd2274: out <= 16'hFFE1;    16'd2275: out <= 16'hFE14;
    16'd2276: out <= 16'hFFAF;    16'd2277: out <= 16'h031B;    16'd2278: out <= 16'hF9A2;    16'd2279: out <= 16'hFE8D;
    16'd2280: out <= 16'h01A5;    16'd2281: out <= 16'h0226;    16'd2282: out <= 16'h0324;    16'd2283: out <= 16'h00B8;
    16'd2284: out <= 16'hFE98;    16'd2285: out <= 16'h056D;    16'd2286: out <= 16'hFDCF;    16'd2287: out <= 16'h027B;
    16'd2288: out <= 16'h0000;    16'd2289: out <= 16'hFD63;    16'd2290: out <= 16'h00A3;    16'd2291: out <= 16'h03D8;
    16'd2292: out <= 16'hFDC2;    16'd2293: out <= 16'h02B3;    16'd2294: out <= 16'h03A4;    16'd2295: out <= 16'h0328;
    16'd2296: out <= 16'hFAB0;    16'd2297: out <= 16'hFD79;    16'd2298: out <= 16'hFD15;    16'd2299: out <= 16'h0534;
    16'd2300: out <= 16'h02A9;    16'd2301: out <= 16'hFB14;    16'd2302: out <= 16'h04BF;    16'd2303: out <= 16'h00D4;
    16'd2304: out <= 16'hFF8B;    16'd2305: out <= 16'h03BA;    16'd2306: out <= 16'h035D;    16'd2307: out <= 16'hF90B;
    16'd2308: out <= 16'h0078;    16'd2309: out <= 16'hFC36;    16'd2310: out <= 16'hFCB8;    16'd2311: out <= 16'hFCD7;
    16'd2312: out <= 16'hFE76;    16'd2313: out <= 16'hFCD1;    16'd2314: out <= 16'hFCFB;    16'd2315: out <= 16'h0209;
    16'd2316: out <= 16'h0007;    16'd2317: out <= 16'h0073;    16'd2318: out <= 16'hFE11;    16'd2319: out <= 16'hFA01;
    16'd2320: out <= 16'h000D;    16'd2321: out <= 16'h0264;    16'd2322: out <= 16'h0135;    16'd2323: out <= 16'hF977;
    16'd2324: out <= 16'hFD6E;    16'd2325: out <= 16'hFBA7;    16'd2326: out <= 16'h0530;    16'd2327: out <= 16'h01A7;
    16'd2328: out <= 16'h01DB;    16'd2329: out <= 16'hFCBF;    16'd2330: out <= 16'h0411;    16'd2331: out <= 16'hFA73;
    16'd2332: out <= 16'hFF81;    16'd2333: out <= 16'h012C;    16'd2334: out <= 16'h00F0;    16'd2335: out <= 16'hFB4F;
    16'd2336: out <= 16'h0919;    16'd2337: out <= 16'hFBD8;    16'd2338: out <= 16'h05CD;    16'd2339: out <= 16'h020F;
    16'd2340: out <= 16'hFF81;    16'd2341: out <= 16'h0198;    16'd2342: out <= 16'h0685;    16'd2343: out <= 16'h04FB;
    16'd2344: out <= 16'h016D;    16'd2345: out <= 16'h03DA;    16'd2346: out <= 16'hFECA;    16'd2347: out <= 16'hFDD6;
    16'd2348: out <= 16'hFA46;    16'd2349: out <= 16'hFD19;    16'd2350: out <= 16'hFDCC;    16'd2351: out <= 16'h0A67;
    16'd2352: out <= 16'h0016;    16'd2353: out <= 16'hFD89;    16'd2354: out <= 16'h06A6;    16'd2355: out <= 16'hFBE8;
    16'd2356: out <= 16'hFE88;    16'd2357: out <= 16'h00DA;    16'd2358: out <= 16'hFA9B;    16'd2359: out <= 16'h074B;
    16'd2360: out <= 16'hFF99;    16'd2361: out <= 16'h05BA;    16'd2362: out <= 16'hFBFE;    16'd2363: out <= 16'hFC58;
    16'd2364: out <= 16'hFB71;    16'd2365: out <= 16'h00FC;    16'd2366: out <= 16'hF8B3;    16'd2367: out <= 16'hFD9A;
    16'd2368: out <= 16'h07DD;    16'd2369: out <= 16'h0655;    16'd2370: out <= 16'h0240;    16'd2371: out <= 16'h032F;
    16'd2372: out <= 16'h08D5;    16'd2373: out <= 16'h0260;    16'd2374: out <= 16'h0025;    16'd2375: out <= 16'h0726;
    16'd2376: out <= 16'h019F;    16'd2377: out <= 16'h03E1;    16'd2378: out <= 16'h0319;    16'd2379: out <= 16'h0520;
    16'd2380: out <= 16'h0809;    16'd2381: out <= 16'h0400;    16'd2382: out <= 16'h0C48;    16'd2383: out <= 16'h000C;
    16'd2384: out <= 16'hFD2C;    16'd2385: out <= 16'h0041;    16'd2386: out <= 16'h01DD;    16'd2387: out <= 16'hFD04;
    16'd2388: out <= 16'hFE0F;    16'd2389: out <= 16'h00A1;    16'd2390: out <= 16'hFA6A;    16'd2391: out <= 16'hFA71;
    16'd2392: out <= 16'h02A7;    16'd2393: out <= 16'hF738;    16'd2394: out <= 16'hFC45;    16'd2395: out <= 16'hFCC7;
    16'd2396: out <= 16'hFA09;    16'd2397: out <= 16'h036D;    16'd2398: out <= 16'hFFA9;    16'd2399: out <= 16'hF6F4;
    16'd2400: out <= 16'hFF75;    16'd2401: out <= 16'h05DB;    16'd2402: out <= 16'hFC38;    16'd2403: out <= 16'h00A7;
    16'd2404: out <= 16'hFE10;    16'd2405: out <= 16'h01C8;    16'd2406: out <= 16'hFBCF;    16'd2407: out <= 16'h048C;
    16'd2408: out <= 16'hFE68;    16'd2409: out <= 16'hFF71;    16'd2410: out <= 16'hFBE2;    16'd2411: out <= 16'hFDC3;
    16'd2412: out <= 16'h05B9;    16'd2413: out <= 16'h0326;    16'd2414: out <= 16'h00E2;    16'd2415: out <= 16'hFDA8;
    16'd2416: out <= 16'h000D;    16'd2417: out <= 16'h0379;    16'd2418: out <= 16'hF9EC;    16'd2419: out <= 16'hFFFB;
    16'd2420: out <= 16'hFEA5;    16'd2421: out <= 16'hF8E6;    16'd2422: out <= 16'hFEB8;    16'd2423: out <= 16'h0224;
    16'd2424: out <= 16'hFD10;    16'd2425: out <= 16'hFC66;    16'd2426: out <= 16'hFDAD;    16'd2427: out <= 16'hFD67;
    16'd2428: out <= 16'h05A1;    16'd2429: out <= 16'h023E;    16'd2430: out <= 16'h02FA;    16'd2431: out <= 16'h06CC;
    16'd2432: out <= 16'hF94C;    16'd2433: out <= 16'h0880;    16'd2434: out <= 16'hFFE2;    16'd2435: out <= 16'hFB78;
    16'd2436: out <= 16'h0590;    16'd2437: out <= 16'h0417;    16'd2438: out <= 16'h07C5;    16'd2439: out <= 16'h0549;
    16'd2440: out <= 16'h058A;    16'd2441: out <= 16'hFD05;    16'd2442: out <= 16'hFD3E;    16'd2443: out <= 16'hFEF5;
    16'd2444: out <= 16'hF719;    16'd2445: out <= 16'h0427;    16'd2446: out <= 16'hFB31;    16'd2447: out <= 16'hFFC5;
    16'd2448: out <= 16'h01E3;    16'd2449: out <= 16'hFE57;    16'd2450: out <= 16'hF847;    16'd2451: out <= 16'hFB93;
    16'd2452: out <= 16'h06FE;    16'd2453: out <= 16'hFC67;    16'd2454: out <= 16'hFB43;    16'd2455: out <= 16'hF90D;
    16'd2456: out <= 16'h05C2;    16'd2457: out <= 16'h020D;    16'd2458: out <= 16'h005C;    16'd2459: out <= 16'hFEC5;
    16'd2460: out <= 16'hFCC1;    16'd2461: out <= 16'hFF8F;    16'd2462: out <= 16'hFFBA;    16'd2463: out <= 16'h004B;
    16'd2464: out <= 16'hFF9D;    16'd2465: out <= 16'h01C9;    16'd2466: out <= 16'hFC6D;    16'd2467: out <= 16'h0344;
    16'd2468: out <= 16'hFD4B;    16'd2469: out <= 16'hFD5E;    16'd2470: out <= 16'h008D;    16'd2471: out <= 16'hFC1F;
    16'd2472: out <= 16'hFF83;    16'd2473: out <= 16'h0731;    16'd2474: out <= 16'h04C1;    16'd2475: out <= 16'h00D0;
    16'd2476: out <= 16'hFFF1;    16'd2477: out <= 16'hFB8F;    16'd2478: out <= 16'hFFAB;    16'd2479: out <= 16'h03C2;
    16'd2480: out <= 16'hFD21;    16'd2481: out <= 16'hFCF1;    16'd2482: out <= 16'hFEBB;    16'd2483: out <= 16'h0164;
    16'd2484: out <= 16'hFD08;    16'd2485: out <= 16'h0181;    16'd2486: out <= 16'hF92D;    16'd2487: out <= 16'h011F;
    16'd2488: out <= 16'h0032;    16'd2489: out <= 16'hFE56;    16'd2490: out <= 16'h01F7;    16'd2491: out <= 16'hFF08;
    16'd2492: out <= 16'h005B;    16'd2493: out <= 16'hFF05;    16'd2494: out <= 16'h013B;    16'd2495: out <= 16'h0362;
    16'd2496: out <= 16'hFB43;    16'd2497: out <= 16'h00C0;    16'd2498: out <= 16'h017E;    16'd2499: out <= 16'h0094;
    16'd2500: out <= 16'hFF4A;    16'd2501: out <= 16'h041D;    16'd2502: out <= 16'hFF76;    16'd2503: out <= 16'hF76F;
    16'd2504: out <= 16'hFCA1;    16'd2505: out <= 16'hFB95;    16'd2506: out <= 16'hFF30;    16'd2507: out <= 16'h0370;
    16'd2508: out <= 16'hFCD2;    16'd2509: out <= 16'h0013;    16'd2510: out <= 16'h025C;    16'd2511: out <= 16'h025E;
    16'd2512: out <= 16'h039D;    16'd2513: out <= 16'h0257;    16'd2514: out <= 16'hFEC4;    16'd2515: out <= 16'h009A;
    16'd2516: out <= 16'h015A;    16'd2517: out <= 16'hFCC2;    16'd2518: out <= 16'h046E;    16'd2519: out <= 16'h00A9;
    16'd2520: out <= 16'h0761;    16'd2521: out <= 16'hFE96;    16'd2522: out <= 16'h0283;    16'd2523: out <= 16'hFCD6;
    16'd2524: out <= 16'hF965;    16'd2525: out <= 16'h018D;    16'd2526: out <= 16'h0036;    16'd2527: out <= 16'h07CF;
    16'd2528: out <= 16'h03A7;    16'd2529: out <= 16'h01EB;    16'd2530: out <= 16'h04B5;    16'd2531: out <= 16'h04E7;
    16'd2532: out <= 16'h0125;    16'd2533: out <= 16'h0460;    16'd2534: out <= 16'h012D;    16'd2535: out <= 16'h0454;
    16'd2536: out <= 16'h01C6;    16'd2537: out <= 16'h023B;    16'd2538: out <= 16'h01CF;    16'd2539: out <= 16'hFF68;
    16'd2540: out <= 16'hFBDF;    16'd2541: out <= 16'h0120;    16'd2542: out <= 16'hFD50;    16'd2543: out <= 16'h01F7;
    16'd2544: out <= 16'h008E;    16'd2545: out <= 16'h03DC;    16'd2546: out <= 16'hFCD0;    16'd2547: out <= 16'h055D;
    16'd2548: out <= 16'h009D;    16'd2549: out <= 16'hFE35;    16'd2550: out <= 16'hFF41;    16'd2551: out <= 16'h078E;
    16'd2552: out <= 16'hFFC7;    16'd2553: out <= 16'h0085;    16'd2554: out <= 16'h018F;    16'd2555: out <= 16'h0853;
    16'd2556: out <= 16'h0234;    16'd2557: out <= 16'hF828;    16'd2558: out <= 16'h0217;    16'd2559: out <= 16'h02CD;
    16'd2560: out <= 16'hF7DA;    16'd2561: out <= 16'hF7E7;    16'd2562: out <= 16'hFE77;    16'd2563: out <= 16'h00BA;
    16'd2564: out <= 16'hFFA2;    16'd2565: out <= 16'hF998;    16'd2566: out <= 16'h02EB;    16'd2567: out <= 16'hF9FC;
    16'd2568: out <= 16'h0163;    16'd2569: out <= 16'h0029;    16'd2570: out <= 16'h093F;    16'd2571: out <= 16'h0447;
    16'd2572: out <= 16'hFFAD;    16'd2573: out <= 16'h0172;    16'd2574: out <= 16'h034E;    16'd2575: out <= 16'h03AD;
    16'd2576: out <= 16'hFC5B;    16'd2577: out <= 16'hFFE5;    16'd2578: out <= 16'h0450;    16'd2579: out <= 16'h02CD;
    16'd2580: out <= 16'hFA47;    16'd2581: out <= 16'hFDC6;    16'd2582: out <= 16'hFF87;    16'd2583: out <= 16'h01E7;
    16'd2584: out <= 16'hFFAE;    16'd2585: out <= 16'hF8B2;    16'd2586: out <= 16'h0A1E;    16'd2587: out <= 16'h00AC;
    16'd2588: out <= 16'h0019;    16'd2589: out <= 16'hFCE4;    16'd2590: out <= 16'h03A4;    16'd2591: out <= 16'hFCEB;
    16'd2592: out <= 16'hFED4;    16'd2593: out <= 16'h036F;    16'd2594: out <= 16'h02E5;    16'd2595: out <= 16'hFDE3;
    16'd2596: out <= 16'h02B7;    16'd2597: out <= 16'hFDC7;    16'd2598: out <= 16'h063D;    16'd2599: out <= 16'h0141;
    16'd2600: out <= 16'h0372;    16'd2601: out <= 16'hFF79;    16'd2602: out <= 16'h0238;    16'd2603: out <= 16'h021F;
    16'd2604: out <= 16'h0673;    16'd2605: out <= 16'hF949;    16'd2606: out <= 16'h0621;    16'd2607: out <= 16'h00E3;
    16'd2608: out <= 16'h003D;    16'd2609: out <= 16'hFA28;    16'd2610: out <= 16'hFFFF;    16'd2611: out <= 16'h01CD;
    16'd2612: out <= 16'h078E;    16'd2613: out <= 16'hFFF8;    16'd2614: out <= 16'hFFFF;    16'd2615: out <= 16'hFD05;
    16'd2616: out <= 16'hFAB6;    16'd2617: out <= 16'h0203;    16'd2618: out <= 16'h0018;    16'd2619: out <= 16'h0549;
    16'd2620: out <= 16'h03A0;    16'd2621: out <= 16'hFCA2;    16'd2622: out <= 16'hFDEE;    16'd2623: out <= 16'h0446;
    16'd2624: out <= 16'hFE5B;    16'd2625: out <= 16'h0547;    16'd2626: out <= 16'hFDAE;    16'd2627: out <= 16'h00C5;
    16'd2628: out <= 16'h0674;    16'd2629: out <= 16'h06D1;    16'd2630: out <= 16'h02B1;    16'd2631: out <= 16'h04BC;
    16'd2632: out <= 16'h0538;    16'd2633: out <= 16'h072B;    16'd2634: out <= 16'h026E;    16'd2635: out <= 16'h04D5;
    16'd2636: out <= 16'h0560;    16'd2637: out <= 16'hFCAF;    16'd2638: out <= 16'h00CD;    16'd2639: out <= 16'h0293;
    16'd2640: out <= 16'hFEC7;    16'd2641: out <= 16'h0623;    16'd2642: out <= 16'h0508;    16'd2643: out <= 16'hFDB5;
    16'd2644: out <= 16'h0704;    16'd2645: out <= 16'hFDD6;    16'd2646: out <= 16'hF786;    16'd2647: out <= 16'h02A2;
    16'd2648: out <= 16'hFE7F;    16'd2649: out <= 16'hF949;    16'd2650: out <= 16'hF6F7;    16'd2651: out <= 16'h00FB;
    16'd2652: out <= 16'h005C;    16'd2653: out <= 16'h0522;    16'd2654: out <= 16'h03BC;    16'd2655: out <= 16'h0853;
    16'd2656: out <= 16'h0094;    16'd2657: out <= 16'h0601;    16'd2658: out <= 16'hFE86;    16'd2659: out <= 16'h00AC;
    16'd2660: out <= 16'h03E9;    16'd2661: out <= 16'hFD02;    16'd2662: out <= 16'hFC05;    16'd2663: out <= 16'hFB72;
    16'd2664: out <= 16'h020E;    16'd2665: out <= 16'hFE56;    16'd2666: out <= 16'hFAFE;    16'd2667: out <= 16'h0012;
    16'd2668: out <= 16'h0222;    16'd2669: out <= 16'h07B4;    16'd2670: out <= 16'h0052;    16'd2671: out <= 16'hFDD4;
    16'd2672: out <= 16'h001A;    16'd2673: out <= 16'hFA67;    16'd2674: out <= 16'h00A6;    16'd2675: out <= 16'h00E2;
    16'd2676: out <= 16'h0492;    16'd2677: out <= 16'h01EA;    16'd2678: out <= 16'hFD3A;    16'd2679: out <= 16'h01FB;
    16'd2680: out <= 16'hFBD7;    16'd2681: out <= 16'hFDBC;    16'd2682: out <= 16'h0337;    16'd2683: out <= 16'h00B5;
    16'd2684: out <= 16'h0480;    16'd2685: out <= 16'hFC29;    16'd2686: out <= 16'hFC3B;    16'd2687: out <= 16'hFBC6;
    16'd2688: out <= 16'h0161;    16'd2689: out <= 16'hFE33;    16'd2690: out <= 16'h03B3;    16'd2691: out <= 16'h0541;
    16'd2692: out <= 16'h0562;    16'd2693: out <= 16'h0836;    16'd2694: out <= 16'h050F;    16'd2695: out <= 16'h0136;
    16'd2696: out <= 16'h0639;    16'd2697: out <= 16'hFB76;    16'd2698: out <= 16'hFE9A;    16'd2699: out <= 16'hFD48;
    16'd2700: out <= 16'h01E5;    16'd2701: out <= 16'hFDC4;    16'd2702: out <= 16'hFAAE;    16'd2703: out <= 16'hFCFB;
    16'd2704: out <= 16'h055B;    16'd2705: out <= 16'h042F;    16'd2706: out <= 16'hFD04;    16'd2707: out <= 16'h0423;
    16'd2708: out <= 16'h026D;    16'd2709: out <= 16'hFE0B;    16'd2710: out <= 16'hFD3A;    16'd2711: out <= 16'h0384;
    16'd2712: out <= 16'hF910;    16'd2713: out <= 16'h0217;    16'd2714: out <= 16'h0567;    16'd2715: out <= 16'hF82C;
    16'd2716: out <= 16'hFA2F;    16'd2717: out <= 16'h005C;    16'd2718: out <= 16'hFE53;    16'd2719: out <= 16'h0281;
    16'd2720: out <= 16'h0450;    16'd2721: out <= 16'h0026;    16'd2722: out <= 16'h05B4;    16'd2723: out <= 16'hFD77;
    16'd2724: out <= 16'h0147;    16'd2725: out <= 16'h0251;    16'd2726: out <= 16'hF9FD;    16'd2727: out <= 16'h0305;
    16'd2728: out <= 16'h088B;    16'd2729: out <= 16'h0348;    16'd2730: out <= 16'hFC20;    16'd2731: out <= 16'hFDEF;
    16'd2732: out <= 16'h012E;    16'd2733: out <= 16'hFB52;    16'd2734: out <= 16'h0AA8;    16'd2735: out <= 16'hFFFE;
    16'd2736: out <= 16'hFE3B;    16'd2737: out <= 16'hFC56;    16'd2738: out <= 16'hFD0F;    16'd2739: out <= 16'hFC3E;
    16'd2740: out <= 16'hF909;    16'd2741: out <= 16'h036B;    16'd2742: out <= 16'h02A2;    16'd2743: out <= 16'h01FF;
    16'd2744: out <= 16'hFEDF;    16'd2745: out <= 16'hFFE1;    16'd2746: out <= 16'hFDD7;    16'd2747: out <= 16'h03C8;
    16'd2748: out <= 16'h0130;    16'd2749: out <= 16'hFD57;    16'd2750: out <= 16'h00E3;    16'd2751: out <= 16'h006C;
    16'd2752: out <= 16'hFC31;    16'd2753: out <= 16'hFEE3;    16'd2754: out <= 16'hFD56;    16'd2755: out <= 16'hFF71;
    16'd2756: out <= 16'h024F;    16'd2757: out <= 16'h05EE;    16'd2758: out <= 16'h00D5;    16'd2759: out <= 16'h008B;
    16'd2760: out <= 16'h00FA;    16'd2761: out <= 16'hFDEA;    16'd2762: out <= 16'h0A5F;    16'd2763: out <= 16'hFCEC;
    16'd2764: out <= 16'hFD98;    16'd2765: out <= 16'h00E7;    16'd2766: out <= 16'h016F;    16'd2767: out <= 16'h00B8;
    16'd2768: out <= 16'h048E;    16'd2769: out <= 16'hFE1F;    16'd2770: out <= 16'hFE2C;    16'd2771: out <= 16'hFFBC;
    16'd2772: out <= 16'hFE4C;    16'd2773: out <= 16'hFC02;    16'd2774: out <= 16'hFEE7;    16'd2775: out <= 16'hFE55;
    16'd2776: out <= 16'h0203;    16'd2777: out <= 16'hF6DF;    16'd2778: out <= 16'hFD00;    16'd2779: out <= 16'hF912;
    16'd2780: out <= 16'h01DF;    16'd2781: out <= 16'h0218;    16'd2782: out <= 16'hFC94;    16'd2783: out <= 16'hFB70;
    16'd2784: out <= 16'hFD1C;    16'd2785: out <= 16'hFDA4;    16'd2786: out <= 16'h024E;    16'd2787: out <= 16'h01A5;
    16'd2788: out <= 16'h01D3;    16'd2789: out <= 16'h0505;    16'd2790: out <= 16'hFC13;    16'd2791: out <= 16'h030D;
    16'd2792: out <= 16'hFD85;    16'd2793: out <= 16'h0119;    16'd2794: out <= 16'h0210;    16'd2795: out <= 16'hFE3E;
    16'd2796: out <= 16'hFF1C;    16'd2797: out <= 16'h017A;    16'd2798: out <= 16'hFC51;    16'd2799: out <= 16'h0142;
    16'd2800: out <= 16'hFEA7;    16'd2801: out <= 16'hFF1F;    16'd2802: out <= 16'h0A7D;    16'd2803: out <= 16'hFA82;
    16'd2804: out <= 16'hFEAC;    16'd2805: out <= 16'hFAD9;    16'd2806: out <= 16'hFD15;    16'd2807: out <= 16'h0072;
    16'd2808: out <= 16'hF8F0;    16'd2809: out <= 16'h07A9;    16'd2810: out <= 16'hFF5E;    16'd2811: out <= 16'hFF6D;
    16'd2812: out <= 16'hFF7C;    16'd2813: out <= 16'hFEFB;    16'd2814: out <= 16'hFDC0;    16'd2815: out <= 16'h026F;
    16'd2816: out <= 16'hF6B6;    16'd2817: out <= 16'h01E0;    16'd2818: out <= 16'h017A;    16'd2819: out <= 16'hFCFA;
    16'd2820: out <= 16'h0198;    16'd2821: out <= 16'hFDB6;    16'd2822: out <= 16'h059E;    16'd2823: out <= 16'hFF10;
    16'd2824: out <= 16'h0206;    16'd2825: out <= 16'h03BF;    16'd2826: out <= 16'hFD9E;    16'd2827: out <= 16'h0010;
    16'd2828: out <= 16'h01B5;    16'd2829: out <= 16'h02CF;    16'd2830: out <= 16'hFEC9;    16'd2831: out <= 16'h004F;
    16'd2832: out <= 16'hFDA7;    16'd2833: out <= 16'hFED8;    16'd2834: out <= 16'hFD2A;    16'd2835: out <= 16'hFE6D;
    16'd2836: out <= 16'h04B7;    16'd2837: out <= 16'h0327;    16'd2838: out <= 16'h000A;    16'd2839: out <= 16'hFC33;
    16'd2840: out <= 16'hFEB4;    16'd2841: out <= 16'hFFDE;    16'd2842: out <= 16'hFD2E;    16'd2843: out <= 16'h048F;
    16'd2844: out <= 16'hFEB3;    16'd2845: out <= 16'hFE36;    16'd2846: out <= 16'h0478;    16'd2847: out <= 16'hFF0C;
    16'd2848: out <= 16'hFAF6;    16'd2849: out <= 16'h0123;    16'd2850: out <= 16'hF849;    16'd2851: out <= 16'hFC75;
    16'd2852: out <= 16'hFAAA;    16'd2853: out <= 16'hFFA2;    16'd2854: out <= 16'hFA2A;    16'd2855: out <= 16'h02C1;
    16'd2856: out <= 16'hF7B9;    16'd2857: out <= 16'h0640;    16'd2858: out <= 16'hFD7A;    16'd2859: out <= 16'hFE45;
    16'd2860: out <= 16'hFFDC;    16'd2861: out <= 16'hFCBC;    16'd2862: out <= 16'h0041;    16'd2863: out <= 16'h0038;
    16'd2864: out <= 16'h04B8;    16'd2865: out <= 16'hFF44;    16'd2866: out <= 16'hF668;    16'd2867: out <= 16'hFE58;
    16'd2868: out <= 16'hF7CF;    16'd2869: out <= 16'h020E;    16'd2870: out <= 16'h029A;    16'd2871: out <= 16'h02EA;
    16'd2872: out <= 16'hFEE6;    16'd2873: out <= 16'hFE8B;    16'd2874: out <= 16'h03BE;    16'd2875: out <= 16'hF6DA;
    16'd2876: out <= 16'hFF48;    16'd2877: out <= 16'h0152;    16'd2878: out <= 16'h0136;    16'd2879: out <= 16'h0521;
    16'd2880: out <= 16'hFD02;    16'd2881: out <= 16'h029D;    16'd2882: out <= 16'h053D;    16'd2883: out <= 16'h03E2;
    16'd2884: out <= 16'h03CC;    16'd2885: out <= 16'h02C3;    16'd2886: out <= 16'hFF90;    16'd2887: out <= 16'h0797;
    16'd2888: out <= 16'h0261;    16'd2889: out <= 16'h016F;    16'd2890: out <= 16'h0020;    16'd2891: out <= 16'h0456;
    16'd2892: out <= 16'h0239;    16'd2893: out <= 16'h064F;    16'd2894: out <= 16'h02C8;    16'd2895: out <= 16'hFF2C;
    16'd2896: out <= 16'h010A;    16'd2897: out <= 16'hF8F5;    16'd2898: out <= 16'h023C;    16'd2899: out <= 16'hFD3D;
    16'd2900: out <= 16'hFE62;    16'd2901: out <= 16'hFA24;    16'd2902: out <= 16'h0011;    16'd2903: out <= 16'h0053;
    16'd2904: out <= 16'hFDA2;    16'd2905: out <= 16'hFBF7;    16'd2906: out <= 16'h0027;    16'd2907: out <= 16'hFD8B;
    16'd2908: out <= 16'hFD14;    16'd2909: out <= 16'hFA9C;    16'd2910: out <= 16'h017C;    16'd2911: out <= 16'h0604;
    16'd2912: out <= 16'h0097;    16'd2913: out <= 16'hFECC;    16'd2914: out <= 16'hFC67;    16'd2915: out <= 16'hFF8C;
    16'd2916: out <= 16'h0041;    16'd2917: out <= 16'h0155;    16'd2918: out <= 16'hFE89;    16'd2919: out <= 16'hFFF4;
    16'd2920: out <= 16'h0685;    16'd2921: out <= 16'hFD10;    16'd2922: out <= 16'hFE05;    16'd2923: out <= 16'h0609;
    16'd2924: out <= 16'h00D6;    16'd2925: out <= 16'hFE25;    16'd2926: out <= 16'hFAF6;    16'd2927: out <= 16'h0349;
    16'd2928: out <= 16'hFE6A;    16'd2929: out <= 16'hFC99;    16'd2930: out <= 16'hFDB5;    16'd2931: out <= 16'h01E3;
    16'd2932: out <= 16'hFE74;    16'd2933: out <= 16'hFCE2;    16'd2934: out <= 16'hFEEF;    16'd2935: out <= 16'hFF34;
    16'd2936: out <= 16'hFEB1;    16'd2937: out <= 16'h0525;    16'd2938: out <= 16'hFE19;    16'd2939: out <= 16'hF84C;
    16'd2940: out <= 16'hFFBF;    16'd2941: out <= 16'h03CC;    16'd2942: out <= 16'hFE3A;    16'd2943: out <= 16'hFE8A;
    16'd2944: out <= 16'h0693;    16'd2945: out <= 16'hF971;    16'd2946: out <= 16'h0490;    16'd2947: out <= 16'h01C2;
    16'd2948: out <= 16'h03AB;    16'd2949: out <= 16'h0604;    16'd2950: out <= 16'h053C;    16'd2951: out <= 16'h017F;
    16'd2952: out <= 16'hFCC3;    16'd2953: out <= 16'h0915;    16'd2954: out <= 16'hFBC0;    16'd2955: out <= 16'hFCAE;
    16'd2956: out <= 16'hFF95;    16'd2957: out <= 16'h01BA;    16'd2958: out <= 16'hFD0E;    16'd2959: out <= 16'hFFD4;
    16'd2960: out <= 16'h04AB;    16'd2961: out <= 16'hF8F1;    16'd2962: out <= 16'hFD3C;    16'd2963: out <= 16'h065E;
    16'd2964: out <= 16'hFD37;    16'd2965: out <= 16'hFCBD;    16'd2966: out <= 16'hF7F6;    16'd2967: out <= 16'h0004;
    16'd2968: out <= 16'hFB73;    16'd2969: out <= 16'h056C;    16'd2970: out <= 16'hFBB9;    16'd2971: out <= 16'h00C5;
    16'd2972: out <= 16'hFF5C;    16'd2973: out <= 16'h09C3;    16'd2974: out <= 16'h01A5;    16'd2975: out <= 16'hFB71;
    16'd2976: out <= 16'hFDFD;    16'd2977: out <= 16'h00AE;    16'd2978: out <= 16'hFC40;    16'd2979: out <= 16'h02F5;
    16'd2980: out <= 16'hFF0A;    16'd2981: out <= 16'h014D;    16'd2982: out <= 16'h01F4;    16'd2983: out <= 16'hFA51;
    16'd2984: out <= 16'hFF22;    16'd2985: out <= 16'hFEA5;    16'd2986: out <= 16'hFB42;    16'd2987: out <= 16'h00A1;
    16'd2988: out <= 16'hFA96;    16'd2989: out <= 16'hFE5C;    16'd2990: out <= 16'h095D;    16'd2991: out <= 16'h015A;
    16'd2992: out <= 16'h006B;    16'd2993: out <= 16'h04F2;    16'd2994: out <= 16'h005C;    16'd2995: out <= 16'h011D;
    16'd2996: out <= 16'h0186;    16'd2997: out <= 16'hF6F3;    16'd2998: out <= 16'h00BC;    16'd2999: out <= 16'h00B2;
    16'd3000: out <= 16'hFD24;    16'd3001: out <= 16'h05E6;    16'd3002: out <= 16'hFB98;    16'd3003: out <= 16'h0136;
    16'd3004: out <= 16'h0340;    16'd3005: out <= 16'h00ED;    16'd3006: out <= 16'h02D0;    16'd3007: out <= 16'h0446;
    16'd3008: out <= 16'h04BF;    16'd3009: out <= 16'hFA9D;    16'd3010: out <= 16'h0121;    16'd3011: out <= 16'hF8B2;
    16'd3012: out <= 16'h00F0;    16'd3013: out <= 16'hFDCE;    16'd3014: out <= 16'h0353;    16'd3015: out <= 16'h0528;
    16'd3016: out <= 16'hFFEC;    16'd3017: out <= 16'hFE65;    16'd3018: out <= 16'hFCC5;    16'd3019: out <= 16'hFE3E;
    16'd3020: out <= 16'hF919;    16'd3021: out <= 16'hFE1B;    16'd3022: out <= 16'h088C;    16'd3023: out <= 16'hF732;
    16'd3024: out <= 16'hFF8E;    16'd3025: out <= 16'h02E3;    16'd3026: out <= 16'hFF19;    16'd3027: out <= 16'hFCD1;
    16'd3028: out <= 16'h03E1;    16'd3029: out <= 16'h02FB;    16'd3030: out <= 16'hFBC3;    16'd3031: out <= 16'hFF25;
    16'd3032: out <= 16'h033C;    16'd3033: out <= 16'hFCB3;    16'd3034: out <= 16'h01E4;    16'd3035: out <= 16'h00A3;
    16'd3036: out <= 16'hFEA5;    16'd3037: out <= 16'hFFE1;    16'd3038: out <= 16'h0265;    16'd3039: out <= 16'h00ED;
    16'd3040: out <= 16'hFD35;    16'd3041: out <= 16'hFCFA;    16'd3042: out <= 16'hFFD7;    16'd3043: out <= 16'hFD56;
    16'd3044: out <= 16'h01A1;    16'd3045: out <= 16'h001D;    16'd3046: out <= 16'hFFE5;    16'd3047: out <= 16'hF9CC;
    16'd3048: out <= 16'hFE84;    16'd3049: out <= 16'h059B;    16'd3050: out <= 16'h059F;    16'd3051: out <= 16'hF967;
    16'd3052: out <= 16'hFD01;    16'd3053: out <= 16'h01BD;    16'd3054: out <= 16'h0193;    16'd3055: out <= 16'hF51B;
    16'd3056: out <= 16'h05D1;    16'd3057: out <= 16'hFF40;    16'd3058: out <= 16'hFD7A;    16'd3059: out <= 16'h0288;
    16'd3060: out <= 16'hFF6F;    16'd3061: out <= 16'hFCE8;    16'd3062: out <= 16'h094A;    16'd3063: out <= 16'hFAD8;
    16'd3064: out <= 16'h025B;    16'd3065: out <= 16'h015F;    16'd3066: out <= 16'h0789;    16'd3067: out <= 16'h02E4;
    16'd3068: out <= 16'h0066;    16'd3069: out <= 16'hFD6C;    16'd3070: out <= 16'hF7BA;    16'd3071: out <= 16'h0621;
    16'd3072: out <= 16'hF6BD;    16'd3073: out <= 16'hFE82;    16'd3074: out <= 16'h0217;    16'd3075: out <= 16'hFF3C;
    16'd3076: out <= 16'h0267;    16'd3077: out <= 16'h04D1;    16'd3078: out <= 16'h00D2;    16'd3079: out <= 16'hF846;
    16'd3080: out <= 16'hFB2A;    16'd3081: out <= 16'hF980;    16'd3082: out <= 16'hFAA8;    16'd3083: out <= 16'hFD10;
    16'd3084: out <= 16'hFFD2;    16'd3085: out <= 16'hFA45;    16'd3086: out <= 16'hFD46;    16'd3087: out <= 16'hFED4;
    16'd3088: out <= 16'hFBA3;    16'd3089: out <= 16'hFA01;    16'd3090: out <= 16'hFE1A;    16'd3091: out <= 16'h044E;
    16'd3092: out <= 16'hFDA5;    16'd3093: out <= 16'h011E;    16'd3094: out <= 16'hF8F9;    16'd3095: out <= 16'h0376;
    16'd3096: out <= 16'hFDE8;    16'd3097: out <= 16'hFFB2;    16'd3098: out <= 16'hFDC1;    16'd3099: out <= 16'h0898;
    16'd3100: out <= 16'hFF34;    16'd3101: out <= 16'hFCD9;    16'd3102: out <= 16'hFA9A;    16'd3103: out <= 16'h0238;
    16'd3104: out <= 16'h0243;    16'd3105: out <= 16'hFD85;    16'd3106: out <= 16'hFED0;    16'd3107: out <= 16'h04D6;
    16'd3108: out <= 16'hFD73;    16'd3109: out <= 16'hFA59;    16'd3110: out <= 16'h05E9;    16'd3111: out <= 16'h048A;
    16'd3112: out <= 16'h0028;    16'd3113: out <= 16'hF62A;    16'd3114: out <= 16'h0420;    16'd3115: out <= 16'h0982;
    16'd3116: out <= 16'hFDFF;    16'd3117: out <= 16'hFC92;    16'd3118: out <= 16'hFBE8;    16'd3119: out <= 16'h0134;
    16'd3120: out <= 16'h01C7;    16'd3121: out <= 16'h0321;    16'd3122: out <= 16'h09AB;    16'd3123: out <= 16'h0545;
    16'd3124: out <= 16'hF958;    16'd3125: out <= 16'h069C;    16'd3126: out <= 16'h010A;    16'd3127: out <= 16'h055C;
    16'd3128: out <= 16'hFE61;    16'd3129: out <= 16'h00DA;    16'd3130: out <= 16'h0101;    16'd3131: out <= 16'hFBD0;
    16'd3132: out <= 16'hFB6D;    16'd3133: out <= 16'h002F;    16'd3134: out <= 16'h0270;    16'd3135: out <= 16'h01E7;
    16'd3136: out <= 16'h085F;    16'd3137: out <= 16'h0280;    16'd3138: out <= 16'hFDDD;    16'd3139: out <= 16'h0456;
    16'd3140: out <= 16'h081C;    16'd3141: out <= 16'h0C3E;    16'd3142: out <= 16'h00F4;    16'd3143: out <= 16'h01F5;
    16'd3144: out <= 16'h0797;    16'd3145: out <= 16'h04C8;    16'd3146: out <= 16'hFF59;    16'd3147: out <= 16'h02BF;
    16'd3148: out <= 16'h0AB4;    16'd3149: out <= 16'hFECC;    16'd3150: out <= 16'h09E3;    16'd3151: out <= 16'hFB56;
    16'd3152: out <= 16'h0206;    16'd3153: out <= 16'h0528;    16'd3154: out <= 16'h0532;    16'd3155: out <= 16'h09F0;
    16'd3156: out <= 16'h0A99;    16'd3157: out <= 16'h0099;    16'd3158: out <= 16'hFD11;    16'd3159: out <= 16'h01C1;
    16'd3160: out <= 16'hFDA2;    16'd3161: out <= 16'h02AB;    16'd3162: out <= 16'h0102;    16'd3163: out <= 16'h02BB;
    16'd3164: out <= 16'h0026;    16'd3165: out <= 16'h0285;    16'd3166: out <= 16'hFE1C;    16'd3167: out <= 16'hF859;
    16'd3168: out <= 16'hF9F9;    16'd3169: out <= 16'hFFBD;    16'd3170: out <= 16'h05B6;    16'd3171: out <= 16'h01E8;
    16'd3172: out <= 16'hFD8B;    16'd3173: out <= 16'hFF3B;    16'd3174: out <= 16'hFFF2;    16'd3175: out <= 16'h06CC;
    16'd3176: out <= 16'hFC26;    16'd3177: out <= 16'hFECF;    16'd3178: out <= 16'h029C;    16'd3179: out <= 16'h0426;
    16'd3180: out <= 16'h03BF;    16'd3181: out <= 16'h0023;    16'd3182: out <= 16'hFEF2;    16'd3183: out <= 16'hFC18;
    16'd3184: out <= 16'h0367;    16'd3185: out <= 16'h0214;    16'd3186: out <= 16'h019A;    16'd3187: out <= 16'hFECB;
    16'd3188: out <= 16'hFD23;    16'd3189: out <= 16'h051A;    16'd3190: out <= 16'h06C3;    16'd3191: out <= 16'h03DA;
    16'd3192: out <= 16'h0193;    16'd3193: out <= 16'h059F;    16'd3194: out <= 16'hFC1A;    16'd3195: out <= 16'hFEF8;
    16'd3196: out <= 16'h0125;    16'd3197: out <= 16'hF852;    16'd3198: out <= 16'hF9DD;    16'd3199: out <= 16'h00DB;
    16'd3200: out <= 16'hFE7C;    16'd3201: out <= 16'h00AA;    16'd3202: out <= 16'hF9EE;    16'd3203: out <= 16'h014C;
    16'd3204: out <= 16'hFD54;    16'd3205: out <= 16'h0526;    16'd3206: out <= 16'h0175;    16'd3207: out <= 16'hFD21;
    16'd3208: out <= 16'hFF9F;    16'd3209: out <= 16'h0383;    16'd3210: out <= 16'hFABD;    16'd3211: out <= 16'hFE93;
    16'd3212: out <= 16'h008A;    16'd3213: out <= 16'h0270;    16'd3214: out <= 16'hFDB8;    16'd3215: out <= 16'h0363;
    16'd3216: out <= 16'h04A7;    16'd3217: out <= 16'h01AC;    16'd3218: out <= 16'hFE54;    16'd3219: out <= 16'hFA21;
    16'd3220: out <= 16'h01B5;    16'd3221: out <= 16'h0420;    16'd3222: out <= 16'h027B;    16'd3223: out <= 16'hFF6A;
    16'd3224: out <= 16'h02C8;    16'd3225: out <= 16'hFBCE;    16'd3226: out <= 16'hFC05;    16'd3227: out <= 16'hFD92;
    16'd3228: out <= 16'h02BF;    16'd3229: out <= 16'hFFD2;    16'd3230: out <= 16'hFF0D;    16'd3231: out <= 16'hFCB4;
    16'd3232: out <= 16'hF56A;    16'd3233: out <= 16'h078A;    16'd3234: out <= 16'hF9B4;    16'd3235: out <= 16'hFEAD;
    16'd3236: out <= 16'hFE60;    16'd3237: out <= 16'hFCD1;    16'd3238: out <= 16'h000B;    16'd3239: out <= 16'hFD53;
    16'd3240: out <= 16'hFEDA;    16'd3241: out <= 16'hF728;    16'd3242: out <= 16'hFDC3;    16'd3243: out <= 16'h0102;
    16'd3244: out <= 16'hF8ED;    16'd3245: out <= 16'hF958;    16'd3246: out <= 16'hFC40;    16'd3247: out <= 16'h0465;
    16'd3248: out <= 16'h0441;    16'd3249: out <= 16'hFE4A;    16'd3250: out <= 16'h04C9;    16'd3251: out <= 16'h031F;
    16'd3252: out <= 16'h000C;    16'd3253: out <= 16'hFE36;    16'd3254: out <= 16'h01AD;    16'd3255: out <= 16'h0497;
    16'd3256: out <= 16'hFC57;    16'd3257: out <= 16'h02B2;    16'd3258: out <= 16'h0358;    16'd3259: out <= 16'h049C;
    16'd3260: out <= 16'hFE1B;    16'd3261: out <= 16'hFE21;    16'd3262: out <= 16'h0269;    16'd3263: out <= 16'hFD9F;
    16'd3264: out <= 16'h00EC;    16'd3265: out <= 16'h0073;    16'd3266: out <= 16'h03BF;    16'd3267: out <= 16'hFF5F;
    16'd3268: out <= 16'h0248;    16'd3269: out <= 16'hFDE5;    16'd3270: out <= 16'h017D;    16'd3271: out <= 16'h02C5;
    16'd3272: out <= 16'hF86A;    16'd3273: out <= 16'hFCA4;    16'd3274: out <= 16'h006B;    16'd3275: out <= 16'h0040;
    16'd3276: out <= 16'hF82D;    16'd3277: out <= 16'hFE4C;    16'd3278: out <= 16'hFF89;    16'd3279: out <= 16'h0476;
    16'd3280: out <= 16'hF815;    16'd3281: out <= 16'h0BBB;    16'd3282: out <= 16'h040C;    16'd3283: out <= 16'h002B;
    16'd3284: out <= 16'hFE0D;    16'd3285: out <= 16'h01E2;    16'd3286: out <= 16'hFBFE;    16'd3287: out <= 16'hFC3D;
    16'd3288: out <= 16'h028E;    16'd3289: out <= 16'h0033;    16'd3290: out <= 16'h01CC;    16'd3291: out <= 16'h0444;
    16'd3292: out <= 16'hFD6D;    16'd3293: out <= 16'h008B;    16'd3294: out <= 16'hFB3B;    16'd3295: out <= 16'h0439;
    16'd3296: out <= 16'h05EF;    16'd3297: out <= 16'hFF56;    16'd3298: out <= 16'h040E;    16'd3299: out <= 16'h01F9;
    16'd3300: out <= 16'h01FA;    16'd3301: out <= 16'hFFCE;    16'd3302: out <= 16'hFBE7;    16'd3303: out <= 16'h047B;
    16'd3304: out <= 16'h0323;    16'd3305: out <= 16'hFDAB;    16'd3306: out <= 16'h0717;    16'd3307: out <= 16'h00CB;
    16'd3308: out <= 16'h0124;    16'd3309: out <= 16'hFE79;    16'd3310: out <= 16'hFA10;    16'd3311: out <= 16'h03C2;
    16'd3312: out <= 16'h014D;    16'd3313: out <= 16'hFFF6;    16'd3314: out <= 16'hFFF4;    16'd3315: out <= 16'h0294;
    16'd3316: out <= 16'hFA07;    16'd3317: out <= 16'h0159;    16'd3318: out <= 16'hFCDA;    16'd3319: out <= 16'h0202;
    16'd3320: out <= 16'h0064;    16'd3321: out <= 16'h00C5;    16'd3322: out <= 16'h0496;    16'd3323: out <= 16'hFBDB;
    16'd3324: out <= 16'h0021;    16'd3325: out <= 16'hF953;    16'd3326: out <= 16'h001D;    16'd3327: out <= 16'hFEB3;
    16'd3328: out <= 16'hFC1D;    16'd3329: out <= 16'hFB26;    16'd3330: out <= 16'h0500;    16'd3331: out <= 16'h0277;
    16'd3332: out <= 16'hFAB4;    16'd3333: out <= 16'h02EA;    16'd3334: out <= 16'h0863;    16'd3335: out <= 16'hFFE0;
    16'd3336: out <= 16'h03E3;    16'd3337: out <= 16'h0095;    16'd3338: out <= 16'hFFCF;    16'd3339: out <= 16'h0761;
    16'd3340: out <= 16'hFB0A;    16'd3341: out <= 16'h028D;    16'd3342: out <= 16'h01B0;    16'd3343: out <= 16'h0365;
    16'd3344: out <= 16'hFB95;    16'd3345: out <= 16'hFF46;    16'd3346: out <= 16'hFB9E;    16'd3347: out <= 16'h0202;
    16'd3348: out <= 16'h07DB;    16'd3349: out <= 16'h02C1;    16'd3350: out <= 16'hFC01;    16'd3351: out <= 16'hFDF0;
    16'd3352: out <= 16'hFFA4;    16'd3353: out <= 16'hFF39;    16'd3354: out <= 16'hFED9;    16'd3355: out <= 16'h0339;
    16'd3356: out <= 16'h00B9;    16'd3357: out <= 16'hF978;    16'd3358: out <= 16'hFE53;    16'd3359: out <= 16'hFBE5;
    16'd3360: out <= 16'hFD94;    16'd3361: out <= 16'h01D7;    16'd3362: out <= 16'h015A;    16'd3363: out <= 16'h02B0;
    16'd3364: out <= 16'hFCE9;    16'd3365: out <= 16'h0029;    16'd3366: out <= 16'h0084;    16'd3367: out <= 16'h0318;
    16'd3368: out <= 16'h04CB;    16'd3369: out <= 16'hFDB1;    16'd3370: out <= 16'hFAAC;    16'd3371: out <= 16'h08DA;
    16'd3372: out <= 16'hF93D;    16'd3373: out <= 16'hFDAC;    16'd3374: out <= 16'hFFF8;    16'd3375: out <= 16'h01E1;
    16'd3376: out <= 16'h0085;    16'd3377: out <= 16'hFA1A;    16'd3378: out <= 16'hFE48;    16'd3379: out <= 16'h023A;
    16'd3380: out <= 16'h030F;    16'd3381: out <= 16'h03FF;    16'd3382: out <= 16'hFDAF;    16'd3383: out <= 16'hFD61;
    16'd3384: out <= 16'h001E;    16'd3385: out <= 16'hF866;    16'd3386: out <= 16'hFC9A;    16'd3387: out <= 16'hFF31;
    16'd3388: out <= 16'h032D;    16'd3389: out <= 16'hFD0B;    16'd3390: out <= 16'h06F9;    16'd3391: out <= 16'h017D;
    16'd3392: out <= 16'h0278;    16'd3393: out <= 16'h02A2;    16'd3394: out <= 16'h01CD;    16'd3395: out <= 16'h0233;
    16'd3396: out <= 16'h06E2;    16'd3397: out <= 16'h0336;    16'd3398: out <= 16'h0465;    16'd3399: out <= 16'h0736;
    16'd3400: out <= 16'h0117;    16'd3401: out <= 16'h029A;    16'd3402: out <= 16'h0665;    16'd3403: out <= 16'hFFE8;
    16'd3404: out <= 16'h0538;    16'd3405: out <= 16'h021B;    16'd3406: out <= 16'h0682;    16'd3407: out <= 16'hFD34;
    16'd3408: out <= 16'h0640;    16'd3409: out <= 16'h0146;    16'd3410: out <= 16'h0657;    16'd3411: out <= 16'h0797;
    16'd3412: out <= 16'h019F;    16'd3413: out <= 16'h072D;    16'd3414: out <= 16'h021C;    16'd3415: out <= 16'h00E4;
    16'd3416: out <= 16'h0615;    16'd3417: out <= 16'h0356;    16'd3418: out <= 16'hFC30;    16'd3419: out <= 16'hFADA;
    16'd3420: out <= 16'h08C1;    16'd3421: out <= 16'h026B;    16'd3422: out <= 16'h01E8;    16'd3423: out <= 16'h0206;
    16'd3424: out <= 16'hFD94;    16'd3425: out <= 16'hF93F;    16'd3426: out <= 16'h0471;    16'd3427: out <= 16'hFEAF;
    16'd3428: out <= 16'h0698;    16'd3429: out <= 16'h048D;    16'd3430: out <= 16'hFF0B;    16'd3431: out <= 16'hFCE3;
    16'd3432: out <= 16'hF941;    16'd3433: out <= 16'h0571;    16'd3434: out <= 16'hFD18;    16'd3435: out <= 16'h037C;
    16'd3436: out <= 16'hF7D5;    16'd3437: out <= 16'hF9E0;    16'd3438: out <= 16'hFC18;    16'd3439: out <= 16'hFD72;
    16'd3440: out <= 16'h04F1;    16'd3441: out <= 16'hFC1B;    16'd3442: out <= 16'hFF9D;    16'd3443: out <= 16'h0469;
    16'd3444: out <= 16'h00AA;    16'd3445: out <= 16'h0114;    16'd3446: out <= 16'hFE38;    16'd3447: out <= 16'h0202;
    16'd3448: out <= 16'hFE0C;    16'd3449: out <= 16'h0043;    16'd3450: out <= 16'hFFAB;    16'd3451: out <= 16'hFE90;
    16'd3452: out <= 16'hFFB6;    16'd3453: out <= 16'h0095;    16'd3454: out <= 16'hFE6C;    16'd3455: out <= 16'h039D;
    16'd3456: out <= 16'h016A;    16'd3457: out <= 16'hFFF0;    16'd3458: out <= 16'h014A;    16'd3459: out <= 16'hFE39;
    16'd3460: out <= 16'hFC23;    16'd3461: out <= 16'hFBF5;    16'd3462: out <= 16'h05C4;    16'd3463: out <= 16'hF902;
    16'd3464: out <= 16'hFED0;    16'd3465: out <= 16'h0036;    16'd3466: out <= 16'h0A7B;    16'd3467: out <= 16'h05CD;
    16'd3468: out <= 16'h072B;    16'd3469: out <= 16'h023A;    16'd3470: out <= 16'hF92B;    16'd3471: out <= 16'h0259;
    16'd3472: out <= 16'h061A;    16'd3473: out <= 16'h034F;    16'd3474: out <= 16'hFE0B;    16'd3475: out <= 16'h02C5;
    16'd3476: out <= 16'h002C;    16'd3477: out <= 16'h018D;    16'd3478: out <= 16'h0394;    16'd3479: out <= 16'hF966;
    16'd3480: out <= 16'hF824;    16'd3481: out <= 16'hFFFD;    16'd3482: out <= 16'hFD4C;    16'd3483: out <= 16'h00B6;
    16'd3484: out <= 16'h0148;    16'd3485: out <= 16'h043B;    16'd3486: out <= 16'hFCD0;    16'd3487: out <= 16'h021C;
    16'd3488: out <= 16'hFE83;    16'd3489: out <= 16'h0409;    16'd3490: out <= 16'h042E;    16'd3491: out <= 16'hFE13;
    16'd3492: out <= 16'hFB78;    16'd3493: out <= 16'h0275;    16'd3494: out <= 16'h0284;    16'd3495: out <= 16'hFE15;
    16'd3496: out <= 16'h05BA;    16'd3497: out <= 16'hFF63;    16'd3498: out <= 16'h00D6;    16'd3499: out <= 16'h00A5;
    16'd3500: out <= 16'h06C1;    16'd3501: out <= 16'h03EF;    16'd3502: out <= 16'h03CA;    16'd3503: out <= 16'hFBEB;
    16'd3504: out <= 16'hFCDA;    16'd3505: out <= 16'h0045;    16'd3506: out <= 16'h00BE;    16'd3507: out <= 16'hFFC7;
    16'd3508: out <= 16'hFD18;    16'd3509: out <= 16'h06E8;    16'd3510: out <= 16'h056B;    16'd3511: out <= 16'h03D1;
    16'd3512: out <= 16'hFCB5;    16'd3513: out <= 16'h00D7;    16'd3514: out <= 16'h00A8;    16'd3515: out <= 16'hFCCD;
    16'd3516: out <= 16'hFAE5;    16'd3517: out <= 16'hFCDB;    16'd3518: out <= 16'hFEFB;    16'd3519: out <= 16'h0212;
    16'd3520: out <= 16'hFABA;    16'd3521: out <= 16'h0420;    16'd3522: out <= 16'h00F6;    16'd3523: out <= 16'h019B;
    16'd3524: out <= 16'hFBB6;    16'd3525: out <= 16'h08DA;    16'd3526: out <= 16'hFCB2;    16'd3527: out <= 16'h03D2;
    16'd3528: out <= 16'h03C4;    16'd3529: out <= 16'h0055;    16'd3530: out <= 16'h031F;    16'd3531: out <= 16'hFF27;
    16'd3532: out <= 16'hFE9B;    16'd3533: out <= 16'h0084;    16'd3534: out <= 16'h03DF;    16'd3535: out <= 16'h0118;
    16'd3536: out <= 16'hFCDE;    16'd3537: out <= 16'h0631;    16'd3538: out <= 16'h0225;    16'd3539: out <= 16'hFE51;
    16'd3540: out <= 16'hFC6B;    16'd3541: out <= 16'h021C;    16'd3542: out <= 16'hFCB3;    16'd3543: out <= 16'h0206;
    16'd3544: out <= 16'h083A;    16'd3545: out <= 16'hFE3B;    16'd3546: out <= 16'h0398;    16'd3547: out <= 16'hFDD9;
    16'd3548: out <= 16'hFFCB;    16'd3549: out <= 16'hFBE9;    16'd3550: out <= 16'hF3DD;    16'd3551: out <= 16'h0014;
    16'd3552: out <= 16'hFF35;    16'd3553: out <= 16'hFF6E;    16'd3554: out <= 16'hFF37;    16'd3555: out <= 16'hFDCB;
    16'd3556: out <= 16'h02D2;    16'd3557: out <= 16'hFF2E;    16'd3558: out <= 16'hFD14;    16'd3559: out <= 16'h0117;
    16'd3560: out <= 16'hFCF1;    16'd3561: out <= 16'hFFEC;    16'd3562: out <= 16'hFFC6;    16'd3563: out <= 16'hFE12;
    16'd3564: out <= 16'hFE0E;    16'd3565: out <= 16'h0760;    16'd3566: out <= 16'h0024;    16'd3567: out <= 16'hFCB5;
    16'd3568: out <= 16'hFF7F;    16'd3569: out <= 16'h0622;    16'd3570: out <= 16'hFBBC;    16'd3571: out <= 16'hFD5C;
    16'd3572: out <= 16'h0018;    16'd3573: out <= 16'h02BB;    16'd3574: out <= 16'h011A;    16'd3575: out <= 16'h031D;
    16'd3576: out <= 16'h0AEB;    16'd3577: out <= 16'h0707;    16'd3578: out <= 16'hFBEB;    16'd3579: out <= 16'h06E8;
    16'd3580: out <= 16'hFF51;    16'd3581: out <= 16'h0160;    16'd3582: out <= 16'h00E4;    16'd3583: out <= 16'h0044;
    16'd3584: out <= 16'hFB6B;    16'd3585: out <= 16'h064F;    16'd3586: out <= 16'hF81D;    16'd3587: out <= 16'h0989;
    16'd3588: out <= 16'hFF0B;    16'd3589: out <= 16'hFF23;    16'd3590: out <= 16'hFF78;    16'd3591: out <= 16'h04CD;
    16'd3592: out <= 16'h0705;    16'd3593: out <= 16'h08FF;    16'd3594: out <= 16'h0400;    16'd3595: out <= 16'hFA0C;
    16'd3596: out <= 16'h0225;    16'd3597: out <= 16'h00FC;    16'd3598: out <= 16'hFE19;    16'd3599: out <= 16'h02FA;
    16'd3600: out <= 16'hFAF1;    16'd3601: out <= 16'h011F;    16'd3602: out <= 16'h0517;    16'd3603: out <= 16'h0342;
    16'd3604: out <= 16'h00B1;    16'd3605: out <= 16'h0197;    16'd3606: out <= 16'h0369;    16'd3607: out <= 16'h0427;
    16'd3608: out <= 16'h032B;    16'd3609: out <= 16'h03BF;    16'd3610: out <= 16'hF9C7;    16'd3611: out <= 16'hFBD6;
    16'd3612: out <= 16'hFCD3;    16'd3613: out <= 16'hFFDE;    16'd3614: out <= 16'h02FE;    16'd3615: out <= 16'h00FD;
    16'd3616: out <= 16'h01A3;    16'd3617: out <= 16'hF832;    16'd3618: out <= 16'hFD52;    16'd3619: out <= 16'hFFA2;
    16'd3620: out <= 16'hFD24;    16'd3621: out <= 16'hFF28;    16'd3622: out <= 16'hFC68;    16'd3623: out <= 16'h0134;
    16'd3624: out <= 16'hFE17;    16'd3625: out <= 16'h015C;    16'd3626: out <= 16'hFF67;    16'd3627: out <= 16'h0205;
    16'd3628: out <= 16'h016C;    16'd3629: out <= 16'hFACA;    16'd3630: out <= 16'h0591;    16'd3631: out <= 16'h0643;
    16'd3632: out <= 16'h08F1;    16'd3633: out <= 16'hFD03;    16'd3634: out <= 16'h0166;    16'd3635: out <= 16'h03D9;
    16'd3636: out <= 16'hFC77;    16'd3637: out <= 16'hFBD9;    16'd3638: out <= 16'h0031;    16'd3639: out <= 16'h0403;
    16'd3640: out <= 16'hFBED;    16'd3641: out <= 16'hF76A;    16'd3642: out <= 16'h032A;    16'd3643: out <= 16'h04E7;
    16'd3644: out <= 16'hFE46;    16'd3645: out <= 16'h01FD;    16'd3646: out <= 16'h0DA4;    16'd3647: out <= 16'hFEE1;
    16'd3648: out <= 16'hFFF2;    16'd3649: out <= 16'h0741;    16'd3650: out <= 16'hFE8F;    16'd3651: out <= 16'h0607;
    16'd3652: out <= 16'hFA96;    16'd3653: out <= 16'h069C;    16'd3654: out <= 16'h0E73;    16'd3655: out <= 16'h0060;
    16'd3656: out <= 16'h0177;    16'd3657: out <= 16'h043A;    16'd3658: out <= 16'h056E;    16'd3659: out <= 16'h0418;
    16'd3660: out <= 16'h06B2;    16'd3661: out <= 16'hFC56;    16'd3662: out <= 16'h02CD;    16'd3663: out <= 16'h06F8;
    16'd3664: out <= 16'h087D;    16'd3665: out <= 16'h0355;    16'd3666: out <= 16'h0C0B;    16'd3667: out <= 16'hF9C8;
    16'd3668: out <= 16'h035A;    16'd3669: out <= 16'hFDC5;    16'd3670: out <= 16'h08F7;    16'd3671: out <= 16'h0698;
    16'd3672: out <= 16'h0557;    16'd3673: out <= 16'h04E8;    16'd3674: out <= 16'h0066;    16'd3675: out <= 16'h0289;
    16'd3676: out <= 16'hFFD6;    16'd3677: out <= 16'h0555;    16'd3678: out <= 16'h055B;    16'd3679: out <= 16'hFB4C;
    16'd3680: out <= 16'hFC91;    16'd3681: out <= 16'hFE5E;    16'd3682: out <= 16'h0431;    16'd3683: out <= 16'hFBFE;
    16'd3684: out <= 16'hFE83;    16'd3685: out <= 16'h0802;    16'd3686: out <= 16'h028A;    16'd3687: out <= 16'hF8D7;
    16'd3688: out <= 16'h013F;    16'd3689: out <= 16'h077C;    16'd3690: out <= 16'h039A;    16'd3691: out <= 16'hFD4C;
    16'd3692: out <= 16'h0036;    16'd3693: out <= 16'hFD3B;    16'd3694: out <= 16'h005A;    16'd3695: out <= 16'h01D5;
    16'd3696: out <= 16'hFB42;    16'd3697: out <= 16'h059E;    16'd3698: out <= 16'h0554;    16'd3699: out <= 16'h0179;
    16'd3700: out <= 16'hFBC2;    16'd3701: out <= 16'hFE99;    16'd3702: out <= 16'h09C4;    16'd3703: out <= 16'h09C5;
    16'd3704: out <= 16'hFF9A;    16'd3705: out <= 16'hFB3C;    16'd3706: out <= 16'hFBBF;    16'd3707: out <= 16'hFEBB;
    16'd3708: out <= 16'hF543;    16'd3709: out <= 16'hFC16;    16'd3710: out <= 16'hF722;    16'd3711: out <= 16'h0080;
    16'd3712: out <= 16'hFEBE;    16'd3713: out <= 16'h043A;    16'd3714: out <= 16'h0117;    16'd3715: out <= 16'hFCD3;
    16'd3716: out <= 16'h0123;    16'd3717: out <= 16'h0036;    16'd3718: out <= 16'hFCF8;    16'd3719: out <= 16'h04E1;
    16'd3720: out <= 16'hFF4F;    16'd3721: out <= 16'hFDA9;    16'd3722: out <= 16'hFCE5;    16'd3723: out <= 16'h00D3;
    16'd3724: out <= 16'hFE9E;    16'd3725: out <= 16'h0678;    16'd3726: out <= 16'h0447;    16'd3727: out <= 16'h0292;
    16'd3728: out <= 16'hFFE1;    16'd3729: out <= 16'h027D;    16'd3730: out <= 16'hFA8C;    16'd3731: out <= 16'hFE46;
    16'd3732: out <= 16'h0385;    16'd3733: out <= 16'h0457;    16'd3734: out <= 16'hFB26;    16'd3735: out <= 16'hFF35;
    16'd3736: out <= 16'h0177;    16'd3737: out <= 16'h0184;    16'd3738: out <= 16'h0064;    16'd3739: out <= 16'hFD88;
    16'd3740: out <= 16'hFBBE;    16'd3741: out <= 16'hFCEA;    16'd3742: out <= 16'hFC44;    16'd3743: out <= 16'hFB5A;
    16'd3744: out <= 16'h034A;    16'd3745: out <= 16'hFEB4;    16'd3746: out <= 16'h0009;    16'd3747: out <= 16'h0250;
    16'd3748: out <= 16'hFAC3;    16'd3749: out <= 16'h0560;    16'd3750: out <= 16'hFB47;    16'd3751: out <= 16'h05DE;
    16'd3752: out <= 16'h0232;    16'd3753: out <= 16'hFEA8;    16'd3754: out <= 16'hF93E;    16'd3755: out <= 16'h01C7;
    16'd3756: out <= 16'h021A;    16'd3757: out <= 16'h02F1;    16'd3758: out <= 16'hFE34;    16'd3759: out <= 16'h0416;
    16'd3760: out <= 16'hFF44;    16'd3761: out <= 16'hFEC6;    16'd3762: out <= 16'h042F;    16'd3763: out <= 16'hFA66;
    16'd3764: out <= 16'h038B;    16'd3765: out <= 16'h037A;    16'd3766: out <= 16'hF6FC;    16'd3767: out <= 16'h0167;
    16'd3768: out <= 16'h0019;    16'd3769: out <= 16'h0408;    16'd3770: out <= 16'hF703;    16'd3771: out <= 16'h03C4;
    16'd3772: out <= 16'hFB10;    16'd3773: out <= 16'hFC31;    16'd3774: out <= 16'h00A0;    16'd3775: out <= 16'h03B9;
    16'd3776: out <= 16'h083D;    16'd3777: out <= 16'h038A;    16'd3778: out <= 16'h0106;    16'd3779: out <= 16'hFA0B;
    16'd3780: out <= 16'h04F3;    16'd3781: out <= 16'h000C;    16'd3782: out <= 16'hFEE8;    16'd3783: out <= 16'hFD73;
    16'd3784: out <= 16'h0243;    16'd3785: out <= 16'h02E5;    16'd3786: out <= 16'h0257;    16'd3787: out <= 16'hFE8C;
    16'd3788: out <= 16'hFFCA;    16'd3789: out <= 16'h0002;    16'd3790: out <= 16'hFA87;    16'd3791: out <= 16'h051C;
    16'd3792: out <= 16'hFFD0;    16'd3793: out <= 16'hFF48;    16'd3794: out <= 16'hFDDF;    16'd3795: out <= 16'hFE02;
    16'd3796: out <= 16'hFFA8;    16'd3797: out <= 16'hFF75;    16'd3798: out <= 16'h0146;    16'd3799: out <= 16'hFBAA;
    16'd3800: out <= 16'h0187;    16'd3801: out <= 16'h0370;    16'd3802: out <= 16'hFE29;    16'd3803: out <= 16'hF958;
    16'd3804: out <= 16'h005C;    16'd3805: out <= 16'h03FC;    16'd3806: out <= 16'hF800;    16'd3807: out <= 16'h0101;
    16'd3808: out <= 16'hFDD0;    16'd3809: out <= 16'hFF3C;    16'd3810: out <= 16'hFDB2;    16'd3811: out <= 16'h04B4;
    16'd3812: out <= 16'h074E;    16'd3813: out <= 16'hFF64;    16'd3814: out <= 16'h00CF;    16'd3815: out <= 16'hF887;
    16'd3816: out <= 16'hFFBF;    16'd3817: out <= 16'h0085;    16'd3818: out <= 16'h006E;    16'd3819: out <= 16'hFFEE;
    16'd3820: out <= 16'h02B4;    16'd3821: out <= 16'hFE59;    16'd3822: out <= 16'h0451;    16'd3823: out <= 16'h011B;
    16'd3824: out <= 16'h0697;    16'd3825: out <= 16'h0AA8;    16'd3826: out <= 16'h011A;    16'd3827: out <= 16'hFFDD;
    16'd3828: out <= 16'h047C;    16'd3829: out <= 16'hFEF0;    16'd3830: out <= 16'h0106;    16'd3831: out <= 16'h020D;
    16'd3832: out <= 16'h0440;    16'd3833: out <= 16'h04A4;    16'd3834: out <= 16'h01C0;    16'd3835: out <= 16'h06F1;
    16'd3836: out <= 16'h038E;    16'd3837: out <= 16'h046B;    16'd3838: out <= 16'h07D6;    16'd3839: out <= 16'hFF9C;
    16'd3840: out <= 16'h03A1;    16'd3841: out <= 16'h06A0;    16'd3842: out <= 16'h0B1B;    16'd3843: out <= 16'hFDE3;
    16'd3844: out <= 16'h0043;    16'd3845: out <= 16'h00EB;    16'd3846: out <= 16'h0638;    16'd3847: out <= 16'hFEFE;
    16'd3848: out <= 16'h0161;    16'd3849: out <= 16'hFF67;    16'd3850: out <= 16'hFF71;    16'd3851: out <= 16'h0264;
    16'd3852: out <= 16'h063F;    16'd3853: out <= 16'h03C6;    16'd3854: out <= 16'h0246;    16'd3855: out <= 16'h05FF;
    16'd3856: out <= 16'hF9FF;    16'd3857: out <= 16'h021C;    16'd3858: out <= 16'h013A;    16'd3859: out <= 16'h0687;
    16'd3860: out <= 16'h04A5;    16'd3861: out <= 16'hFF6E;    16'd3862: out <= 16'h0568;    16'd3863: out <= 16'hFE8B;
    16'd3864: out <= 16'hFA56;    16'd3865: out <= 16'h051E;    16'd3866: out <= 16'h051F;    16'd3867: out <= 16'hF4D7;
    16'd3868: out <= 16'hFF0C;    16'd3869: out <= 16'h009C;    16'd3870: out <= 16'hFA3A;    16'd3871: out <= 16'h01B4;
    16'd3872: out <= 16'hFEE1;    16'd3873: out <= 16'hFFB7;    16'd3874: out <= 16'hFD6B;    16'd3875: out <= 16'hFE0E;
    16'd3876: out <= 16'h03C4;    16'd3877: out <= 16'hFC51;    16'd3878: out <= 16'hFE58;    16'd3879: out <= 16'hFE3C;
    16'd3880: out <= 16'h008D;    16'd3881: out <= 16'h082B;    16'd3882: out <= 16'h0091;    16'd3883: out <= 16'hFA7A;
    16'd3884: out <= 16'hFBD2;    16'd3885: out <= 16'h03FA;    16'd3886: out <= 16'hFD7B;    16'd3887: out <= 16'h030B;
    16'd3888: out <= 16'hFA07;    16'd3889: out <= 16'hFF88;    16'd3890: out <= 16'h0276;    16'd3891: out <= 16'h022F;
    16'd3892: out <= 16'h0120;    16'd3893: out <= 16'h0B2E;    16'd3894: out <= 16'h00F4;    16'd3895: out <= 16'hFB73;
    16'd3896: out <= 16'h00E8;    16'd3897: out <= 16'h02E5;    16'd3898: out <= 16'hFFC8;    16'd3899: out <= 16'h037E;
    16'd3900: out <= 16'h038B;    16'd3901: out <= 16'h0485;    16'd3902: out <= 16'h0943;    16'd3903: out <= 16'h07CD;
    16'd3904: out <= 16'h0454;    16'd3905: out <= 16'h05EC;    16'd3906: out <= 16'h017D;    16'd3907: out <= 16'h0355;
    16'd3908: out <= 16'h09C1;    16'd3909: out <= 16'h09F8;    16'd3910: out <= 16'h022B;    16'd3911: out <= 16'h02EE;
    16'd3912: out <= 16'h0351;    16'd3913: out <= 16'h0071;    16'd3914: out <= 16'h085E;    16'd3915: out <= 16'hFFD7;
    16'd3916: out <= 16'h02EE;    16'd3917: out <= 16'h065E;    16'd3918: out <= 16'h01F5;    16'd3919: out <= 16'h03EF;
    16'd3920: out <= 16'h023D;    16'd3921: out <= 16'h00DA;    16'd3922: out <= 16'h0821;    16'd3923: out <= 16'h058B;
    16'd3924: out <= 16'h008A;    16'd3925: out <= 16'h0865;    16'd3926: out <= 16'h038A;    16'd3927: out <= 16'h021D;
    16'd3928: out <= 16'h04D5;    16'd3929: out <= 16'h033A;    16'd3930: out <= 16'h0444;    16'd3931: out <= 16'hFCC4;
    16'd3932: out <= 16'h08BE;    16'd3933: out <= 16'h0114;    16'd3934: out <= 16'h0B3F;    16'd3935: out <= 16'h0808;
    16'd3936: out <= 16'h0252;    16'd3937: out <= 16'h0254;    16'd3938: out <= 16'h060A;    16'd3939: out <= 16'hFBE8;
    16'd3940: out <= 16'hFE53;    16'd3941: out <= 16'hFD9C;    16'd3942: out <= 16'h02CE;    16'd3943: out <= 16'h04E7;
    16'd3944: out <= 16'h0163;    16'd3945: out <= 16'h03C4;    16'd3946: out <= 16'hFD0B;    16'd3947: out <= 16'h0007;
    16'd3948: out <= 16'hFB57;    16'd3949: out <= 16'hF9DA;    16'd3950: out <= 16'hFF9E;    16'd3951: out <= 16'h0193;
    16'd3952: out <= 16'hFBED;    16'd3953: out <= 16'h06E8;    16'd3954: out <= 16'h05EF;    16'd3955: out <= 16'hFE87;
    16'd3956: out <= 16'hFC51;    16'd3957: out <= 16'h05BC;    16'd3958: out <= 16'h0196;    16'd3959: out <= 16'hFFA5;
    16'd3960: out <= 16'h0386;    16'd3961: out <= 16'h06E8;    16'd3962: out <= 16'h0548;    16'd3963: out <= 16'h076C;
    16'd3964: out <= 16'hFADD;    16'd3965: out <= 16'h06D9;    16'd3966: out <= 16'h02CF;    16'd3967: out <= 16'h04DE;
    16'd3968: out <= 16'h000D;    16'd3969: out <= 16'hFDF2;    16'd3970: out <= 16'h024F;    16'd3971: out <= 16'hFC2B;
    16'd3972: out <= 16'h049E;    16'd3973: out <= 16'h05AC;    16'd3974: out <= 16'h03EB;    16'd3975: out <= 16'h074F;
    16'd3976: out <= 16'hFFFA;    16'd3977: out <= 16'h0AFD;    16'd3978: out <= 16'h0292;    16'd3979: out <= 16'h0705;
    16'd3980: out <= 16'h0260;    16'd3981: out <= 16'hF90B;    16'd3982: out <= 16'hF8A0;    16'd3983: out <= 16'h0629;
    16'd3984: out <= 16'h0433;    16'd3985: out <= 16'h0149;    16'd3986: out <= 16'h0027;    16'd3987: out <= 16'h002E;
    16'd3988: out <= 16'h02F6;    16'd3989: out <= 16'h06AC;    16'd3990: out <= 16'hFC4D;    16'd3991: out <= 16'hFDF2;
    16'd3992: out <= 16'hF7BF;    16'd3993: out <= 16'h0305;    16'd3994: out <= 16'h0218;    16'd3995: out <= 16'hFFA3;
    16'd3996: out <= 16'hFABF;    16'd3997: out <= 16'h0091;    16'd3998: out <= 16'hF96B;    16'd3999: out <= 16'hFE3E;
    16'd4000: out <= 16'hFC81;    16'd4001: out <= 16'h0573;    16'd4002: out <= 16'hFF45;    16'd4003: out <= 16'hFF35;
    16'd4004: out <= 16'h02CC;    16'd4005: out <= 16'hFFEE;    16'd4006: out <= 16'h02CD;    16'd4007: out <= 16'hFBE1;
    16'd4008: out <= 16'hFEE7;    16'd4009: out <= 16'h04CA;    16'd4010: out <= 16'h06E7;    16'd4011: out <= 16'h0270;
    16'd4012: out <= 16'h0349;    16'd4013: out <= 16'h047E;    16'd4014: out <= 16'h0495;    16'd4015: out <= 16'hFC84;
    16'd4016: out <= 16'h02AC;    16'd4017: out <= 16'h000F;    16'd4018: out <= 16'h00CC;    16'd4019: out <= 16'hFEDC;
    16'd4020: out <= 16'h0447;    16'd4021: out <= 16'h04F1;    16'd4022: out <= 16'h0057;    16'd4023: out <= 16'h016B;
    16'd4024: out <= 16'h002B;    16'd4025: out <= 16'h033E;    16'd4026: out <= 16'h0408;    16'd4027: out <= 16'h0162;
    16'd4028: out <= 16'h09B1;    16'd4029: out <= 16'h0153;    16'd4030: out <= 16'hFD70;    16'd4031: out <= 16'h0191;
    16'd4032: out <= 16'h0676;    16'd4033: out <= 16'h0267;    16'd4034: out <= 16'hFA56;    16'd4035: out <= 16'h03B5;
    16'd4036: out <= 16'h029F;    16'd4037: out <= 16'h0481;    16'd4038: out <= 16'hF95F;    16'd4039: out <= 16'h06C2;
    16'd4040: out <= 16'hFEDD;    16'd4041: out <= 16'hFEAF;    16'd4042: out <= 16'hFFBE;    16'd4043: out <= 16'hFF6F;
    16'd4044: out <= 16'h017D;    16'd4045: out <= 16'h00F3;    16'd4046: out <= 16'h0AF1;    16'd4047: out <= 16'hF9DA;
    16'd4048: out <= 16'hFBA1;    16'd4049: out <= 16'h0449;    16'd4050: out <= 16'h0370;    16'd4051: out <= 16'h03E2;
    16'd4052: out <= 16'h03A0;    16'd4053: out <= 16'hFE11;    16'd4054: out <= 16'hF822;    16'd4055: out <= 16'h0039;
    16'd4056: out <= 16'hFD4E;    16'd4057: out <= 16'hFFE4;    16'd4058: out <= 16'hFF08;    16'd4059: out <= 16'h00FF;
    16'd4060: out <= 16'h001F;    16'd4061: out <= 16'hFF3E;    16'd4062: out <= 16'h0112;    16'd4063: out <= 16'h0358;
    16'd4064: out <= 16'hFF9C;    16'd4065: out <= 16'hFE41;    16'd4066: out <= 16'hFC98;    16'd4067: out <= 16'h0200;
    16'd4068: out <= 16'hFDF7;    16'd4069: out <= 16'hFD2C;    16'd4070: out <= 16'h047C;    16'd4071: out <= 16'hFEF0;
    16'd4072: out <= 16'h0073;    16'd4073: out <= 16'hFFE4;    16'd4074: out <= 16'hFD0C;    16'd4075: out <= 16'h068A;
    16'd4076: out <= 16'hFFBD;    16'd4077: out <= 16'h0124;    16'd4078: out <= 16'hFCE7;    16'd4079: out <= 16'hF7DA;
    16'd4080: out <= 16'hFA02;    16'd4081: out <= 16'h0293;    16'd4082: out <= 16'hF7D7;    16'd4083: out <= 16'hFF44;
    16'd4084: out <= 16'h05FC;    16'd4085: out <= 16'h02D3;    16'd4086: out <= 16'hF937;    16'd4087: out <= 16'hFBC1;
    16'd4088: out <= 16'h02A5;    16'd4089: out <= 16'hF9C6;    16'd4090: out <= 16'h01C0;    16'd4091: out <= 16'hFCFB;
    16'd4092: out <= 16'h0285;    16'd4093: out <= 16'hFFEC;    16'd4094: out <= 16'hFD54;    16'd4095: out <= 16'hFBF0;
    16'd4096: out <= 16'h0312;    16'd4097: out <= 16'h002B;    16'd4098: out <= 16'hFE57;    16'd4099: out <= 16'h049F;
    16'd4100: out <= 16'hFEB9;    16'd4101: out <= 16'h0236;    16'd4102: out <= 16'hFD41;    16'd4103: out <= 16'h02C2;
    16'd4104: out <= 16'hFC90;    16'd4105: out <= 16'h04BA;    16'd4106: out <= 16'hF8E6;    16'd4107: out <= 16'h01C2;
    16'd4108: out <= 16'h06DD;    16'd4109: out <= 16'hFAF7;    16'd4110: out <= 16'h00B5;    16'd4111: out <= 16'h02CD;
    16'd4112: out <= 16'hFEBA;    16'd4113: out <= 16'hFD8F;    16'd4114: out <= 16'h0734;    16'd4115: out <= 16'h01FB;
    16'd4116: out <= 16'h0441;    16'd4117: out <= 16'h0584;    16'd4118: out <= 16'hFF57;    16'd4119: out <= 16'hFA7F;
    16'd4120: out <= 16'h02C5;    16'd4121: out <= 16'hF95F;    16'd4122: out <= 16'hFD16;    16'd4123: out <= 16'h0A92;
    16'd4124: out <= 16'hFE4F;    16'd4125: out <= 16'hFA64;    16'd4126: out <= 16'hFCA4;    16'd4127: out <= 16'hFDB8;
    16'd4128: out <= 16'h00A6;    16'd4129: out <= 16'hF890;    16'd4130: out <= 16'hFCB1;    16'd4131: out <= 16'h045F;
    16'd4132: out <= 16'hFC41;    16'd4133: out <= 16'h050D;    16'd4134: out <= 16'h0312;    16'd4135: out <= 16'hFD6B;
    16'd4136: out <= 16'h0268;    16'd4137: out <= 16'h0110;    16'd4138: out <= 16'hFB28;    16'd4139: out <= 16'hFAEF;
    16'd4140: out <= 16'hFC7D;    16'd4141: out <= 16'h02A1;    16'd4142: out <= 16'h0695;    16'd4143: out <= 16'hFD37;
    16'd4144: out <= 16'h0552;    16'd4145: out <= 16'h0138;    16'd4146: out <= 16'h08BE;    16'd4147: out <= 16'hFD91;
    16'd4148: out <= 16'h069C;    16'd4149: out <= 16'h05EA;    16'd4150: out <= 16'h0252;    16'd4151: out <= 16'h01AB;
    16'd4152: out <= 16'hF757;    16'd4153: out <= 16'h00B3;    16'd4154: out <= 16'h03D0;    16'd4155: out <= 16'h03EB;
    16'd4156: out <= 16'h0B49;    16'd4157: out <= 16'h06D4;    16'd4158: out <= 16'h07D4;    16'd4159: out <= 16'h07B0;
    16'd4160: out <= 16'h0C1E;    16'd4161: out <= 16'h0093;    16'd4162: out <= 16'h0523;    16'd4163: out <= 16'h06C6;
    16'd4164: out <= 16'h0C81;    16'd4165: out <= 16'h050F;    16'd4166: out <= 16'hFBE8;    16'd4167: out <= 16'h06AB;
    16'd4168: out <= 16'h041A;    16'd4169: out <= 16'h03F8;    16'd4170: out <= 16'h095A;    16'd4171: out <= 16'h0A39;
    16'd4172: out <= 16'h0A30;    16'd4173: out <= 16'h069F;    16'd4174: out <= 16'h04E5;    16'd4175: out <= 16'h046F;
    16'd4176: out <= 16'h02B7;    16'd4177: out <= 16'h02F9;    16'd4178: out <= 16'h035F;    16'd4179: out <= 16'h0A58;
    16'd4180: out <= 16'h00D8;    16'd4181: out <= 16'h05E9;    16'd4182: out <= 16'h01BD;    16'd4183: out <= 16'h0705;
    16'd4184: out <= 16'hFE40;    16'd4185: out <= 16'h02DB;    16'd4186: out <= 16'h0717;    16'd4187: out <= 16'h08B2;
    16'd4188: out <= 16'h05BE;    16'd4189: out <= 16'h0797;    16'd4190: out <= 16'hFFE2;    16'd4191: out <= 16'h0656;
    16'd4192: out <= 16'h00F2;    16'd4193: out <= 16'h01C3;    16'd4194: out <= 16'h0414;    16'd4195: out <= 16'h094B;
    16'd4196: out <= 16'h00E0;    16'd4197: out <= 16'h01BD;    16'd4198: out <= 16'h0147;    16'd4199: out <= 16'h01CB;
    16'd4200: out <= 16'h08D0;    16'd4201: out <= 16'h0232;    16'd4202: out <= 16'h0175;    16'd4203: out <= 16'hFF18;
    16'd4204: out <= 16'h0327;    16'd4205: out <= 16'h038F;    16'd4206: out <= 16'h0756;    16'd4207: out <= 16'hFFCC;
    16'd4208: out <= 16'hFE88;    16'd4209: out <= 16'h01A3;    16'd4210: out <= 16'h0576;    16'd4211: out <= 16'h02EF;
    16'd4212: out <= 16'hFF6C;    16'd4213: out <= 16'h0C4A;    16'd4214: out <= 16'h0CF7;    16'd4215: out <= 16'hFF15;
    16'd4216: out <= 16'h03C3;    16'd4217: out <= 16'h04F0;    16'd4218: out <= 16'hFFA8;    16'd4219: out <= 16'h0873;
    16'd4220: out <= 16'h07C1;    16'd4221: out <= 16'hFEEE;    16'd4222: out <= 16'h0132;    16'd4223: out <= 16'h06AF;
    16'd4224: out <= 16'h09AA;    16'd4225: out <= 16'h04C8;    16'd4226: out <= 16'h0660;    16'd4227: out <= 16'h054E;
    16'd4228: out <= 16'h041C;    16'd4229: out <= 16'h0553;    16'd4230: out <= 16'h0BE1;    16'd4231: out <= 16'hFB59;
    16'd4232: out <= 16'hFE73;    16'd4233: out <= 16'h01ED;    16'd4234: out <= 16'h02A9;    16'd4235: out <= 16'hF9E0;
    16'd4236: out <= 16'h01B9;    16'd4237: out <= 16'hFFB2;    16'd4238: out <= 16'h02F3;    16'd4239: out <= 16'hFD09;
    16'd4240: out <= 16'hFB59;    16'd4241: out <= 16'hFD6B;    16'd4242: out <= 16'hFEA9;    16'd4243: out <= 16'h02C2;
    16'd4244: out <= 16'h0042;    16'd4245: out <= 16'h07CC;    16'd4246: out <= 16'hFF71;    16'd4247: out <= 16'hFE60;
    16'd4248: out <= 16'h00F6;    16'd4249: out <= 16'hFD42;    16'd4250: out <= 16'h00FE;    16'd4251: out <= 16'h0248;
    16'd4252: out <= 16'hFBC1;    16'd4253: out <= 16'hFD53;    16'd4254: out <= 16'h014E;    16'd4255: out <= 16'hFC88;
    16'd4256: out <= 16'hFA71;    16'd4257: out <= 16'h0446;    16'd4258: out <= 16'hFDD6;    16'd4259: out <= 16'hFFBF;
    16'd4260: out <= 16'h02A2;    16'd4261: out <= 16'h0103;    16'd4262: out <= 16'hFD65;    16'd4263: out <= 16'h02AE;
    16'd4264: out <= 16'h057A;    16'd4265: out <= 16'hFF39;    16'd4266: out <= 16'hFFB8;    16'd4267: out <= 16'h046F;
    16'd4268: out <= 16'h0341;    16'd4269: out <= 16'hFE61;    16'd4270: out <= 16'h00DD;    16'd4271: out <= 16'h09A9;
    16'd4272: out <= 16'h0658;    16'd4273: out <= 16'h04BF;    16'd4274: out <= 16'h03ED;    16'd4275: out <= 16'h04BC;
    16'd4276: out <= 16'h0817;    16'd4277: out <= 16'hFCAE;    16'd4278: out <= 16'hF87F;    16'd4279: out <= 16'hFD3C;
    16'd4280: out <= 16'h03E0;    16'd4281: out <= 16'h02B9;    16'd4282: out <= 16'h061B;    16'd4283: out <= 16'h0068;
    16'd4284: out <= 16'h04B4;    16'd4285: out <= 16'hFD7E;    16'd4286: out <= 16'h03FB;    16'd4287: out <= 16'hFFA8;
    16'd4288: out <= 16'hFC4A;    16'd4289: out <= 16'hFB45;    16'd4290: out <= 16'h00DE;    16'd4291: out <= 16'hFB2B;
    16'd4292: out <= 16'hFB8F;    16'd4293: out <= 16'hFC79;    16'd4294: out <= 16'h02A9;    16'd4295: out <= 16'hFE28;
    16'd4296: out <= 16'hFF83;    16'd4297: out <= 16'h0317;    16'd4298: out <= 16'hFFFF;    16'd4299: out <= 16'hFF08;
    16'd4300: out <= 16'hFE7D;    16'd4301: out <= 16'h08FB;    16'd4302: out <= 16'h0680;    16'd4303: out <= 16'h054B;
    16'd4304: out <= 16'h0674;    16'd4305: out <= 16'hF95F;    16'd4306: out <= 16'h02CD;    16'd4307: out <= 16'h02BF;
    16'd4308: out <= 16'h019C;    16'd4309: out <= 16'h0129;    16'd4310: out <= 16'hFEFE;    16'd4311: out <= 16'h0511;
    16'd4312: out <= 16'hFC9B;    16'd4313: out <= 16'h0066;    16'd4314: out <= 16'hFF27;    16'd4315: out <= 16'hFDB5;
    16'd4316: out <= 16'hFF90;    16'd4317: out <= 16'h020F;    16'd4318: out <= 16'h02CF;    16'd4319: out <= 16'hFAFD;
    16'd4320: out <= 16'hFB3E;    16'd4321: out <= 16'hFF0C;    16'd4322: out <= 16'h02E3;    16'd4323: out <= 16'h01D7;
    16'd4324: out <= 16'h0349;    16'd4325: out <= 16'hFF42;    16'd4326: out <= 16'h0114;    16'd4327: out <= 16'hFA35;
    16'd4328: out <= 16'hFDE8;    16'd4329: out <= 16'hFC99;    16'd4330: out <= 16'hFAE6;    16'd4331: out <= 16'hFD11;
    16'd4332: out <= 16'h0575;    16'd4333: out <= 16'hF6B0;    16'd4334: out <= 16'hFD7B;    16'd4335: out <= 16'h0134;
    16'd4336: out <= 16'hFB56;    16'd4337: out <= 16'h0559;    16'd4338: out <= 16'h00A8;    16'd4339: out <= 16'hFF07;
    16'd4340: out <= 16'hFBA9;    16'd4341: out <= 16'h0007;    16'd4342: out <= 16'h0064;    16'd4343: out <= 16'h02ED;
    16'd4344: out <= 16'hFF49;    16'd4345: out <= 16'h0044;    16'd4346: out <= 16'hF60A;    16'd4347: out <= 16'hFD24;
    16'd4348: out <= 16'h0030;    16'd4349: out <= 16'hFEF4;    16'd4350: out <= 16'h05BA;    16'd4351: out <= 16'hFE01;
    16'd4352: out <= 16'h01E7;    16'd4353: out <= 16'hF4A7;    16'd4354: out <= 16'hF91D;    16'd4355: out <= 16'h0320;
    16'd4356: out <= 16'h0275;    16'd4357: out <= 16'hFA6B;    16'd4358: out <= 16'h0434;    16'd4359: out <= 16'h0443;
    16'd4360: out <= 16'h05C9;    16'd4361: out <= 16'h0167;    16'd4362: out <= 16'h002A;    16'd4363: out <= 16'hFB9F;
    16'd4364: out <= 16'h0029;    16'd4365: out <= 16'hFDA7;    16'd4366: out <= 16'h0017;    16'd4367: out <= 16'h0026;
    16'd4368: out <= 16'h044C;    16'd4369: out <= 16'h02DF;    16'd4370: out <= 16'hFD0A;    16'd4371: out <= 16'hF98F;
    16'd4372: out <= 16'h06D0;    16'd4373: out <= 16'hFE67;    16'd4374: out <= 16'hFDCE;    16'd4375: out <= 16'hFCB2;
    16'd4376: out <= 16'hFE2F;    16'd4377: out <= 16'hFFAF;    16'd4378: out <= 16'h0405;    16'd4379: out <= 16'h0389;
    16'd4380: out <= 16'hFEF0;    16'd4381: out <= 16'h0100;    16'd4382: out <= 16'hFB0F;    16'd4383: out <= 16'h0779;
    16'd4384: out <= 16'h0353;    16'd4385: out <= 16'hFAB4;    16'd4386: out <= 16'h0172;    16'd4387: out <= 16'hFB4B;
    16'd4388: out <= 16'hFF5A;    16'd4389: out <= 16'hFA13;    16'd4390: out <= 16'hFC47;    16'd4391: out <= 16'hFB03;
    16'd4392: out <= 16'hF356;    16'd4393: out <= 16'hFE64;    16'd4394: out <= 16'hFF12;    16'd4395: out <= 16'h0218;
    16'd4396: out <= 16'hF9FC;    16'd4397: out <= 16'hFEDB;    16'd4398: out <= 16'h05E4;    16'd4399: out <= 16'h0609;
    16'd4400: out <= 16'h037D;    16'd4401: out <= 16'h01AE;    16'd4402: out <= 16'h00F4;    16'd4403: out <= 16'hFC5A;
    16'd4404: out <= 16'hFFD7;    16'd4405: out <= 16'h039D;    16'd4406: out <= 16'h00AB;    16'd4407: out <= 16'hFD57;
    16'd4408: out <= 16'h0600;    16'd4409: out <= 16'h0280;    16'd4410: out <= 16'h066D;    16'd4411: out <= 16'h06D4;
    16'd4412: out <= 16'h0745;    16'd4413: out <= 16'h0106;    16'd4414: out <= 16'h0484;    16'd4415: out <= 16'hFFB4;
    16'd4416: out <= 16'h0992;    16'd4417: out <= 16'h0432;    16'd4418: out <= 16'h030D;    16'd4419: out <= 16'h031D;
    16'd4420: out <= 16'h07A0;    16'd4421: out <= 16'h06FB;    16'd4422: out <= 16'hFF09;    16'd4423: out <= 16'h0A18;
    16'd4424: out <= 16'h0313;    16'd4425: out <= 16'h08EE;    16'd4426: out <= 16'h013A;    16'd4427: out <= 16'h0454;
    16'd4428: out <= 16'h011E;    16'd4429: out <= 16'h02C8;    16'd4430: out <= 16'h0466;    16'd4431: out <= 16'h0284;
    16'd4432: out <= 16'h0299;    16'd4433: out <= 16'h0094;    16'd4434: out <= 16'h0450;    16'd4435: out <= 16'h0577;
    16'd4436: out <= 16'h06CE;    16'd4437: out <= 16'h00E0;    16'd4438: out <= 16'h00B1;    16'd4439: out <= 16'h02D9;
    16'd4440: out <= 16'h01C4;    16'd4441: out <= 16'h0198;    16'd4442: out <= 16'h079A;    16'd4443: out <= 16'h0BD7;
    16'd4444: out <= 16'h032A;    16'd4445: out <= 16'h055B;    16'd4446: out <= 16'h0630;    16'd4447: out <= 16'hFE10;
    16'd4448: out <= 16'h055C;    16'd4449: out <= 16'h09A9;    16'd4450: out <= 16'hFC89;    16'd4451: out <= 16'h0422;
    16'd4452: out <= 16'h0174;    16'd4453: out <= 16'h0990;    16'd4454: out <= 16'h0891;    16'd4455: out <= 16'h056E;
    16'd4456: out <= 16'h0489;    16'd4457: out <= 16'h0323;    16'd4458: out <= 16'h0D84;    16'd4459: out <= 16'h041A;
    16'd4460: out <= 16'h0204;    16'd4461: out <= 16'h04E9;    16'd4462: out <= 16'hFD9F;    16'd4463: out <= 16'h01CC;
    16'd4464: out <= 16'h06E4;    16'd4465: out <= 16'h076B;    16'd4466: out <= 16'h0026;    16'd4467: out <= 16'h0DAE;
    16'd4468: out <= 16'h03A6;    16'd4469: out <= 16'h0242;    16'd4470: out <= 16'h0547;    16'd4471: out <= 16'h08D6;
    16'd4472: out <= 16'h0295;    16'd4473: out <= 16'hFC1C;    16'd4474: out <= 16'h08DD;    16'd4475: out <= 16'h0012;
    16'd4476: out <= 16'h058F;    16'd4477: out <= 16'h0229;    16'd4478: out <= 16'h05C6;    16'd4479: out <= 16'h0028;
    16'd4480: out <= 16'h0500;    16'd4481: out <= 16'h07E3;    16'd4482: out <= 16'hFF6B;    16'd4483: out <= 16'h04E7;
    16'd4484: out <= 16'hFAD5;    16'd4485: out <= 16'h0A5D;    16'd4486: out <= 16'h0B19;    16'd4487: out <= 16'h0350;
    16'd4488: out <= 16'hFFEC;    16'd4489: out <= 16'h0489;    16'd4490: out <= 16'h036D;    16'd4491: out <= 16'h0691;
    16'd4492: out <= 16'h0926;    16'd4493: out <= 16'h02D0;    16'd4494: out <= 16'h07BD;    16'd4495: out <= 16'h033D;
    16'd4496: out <= 16'h08C0;    16'd4497: out <= 16'h00F3;    16'd4498: out <= 16'hFF1C;    16'd4499: out <= 16'h017A;
    16'd4500: out <= 16'h01D6;    16'd4501: out <= 16'h037C;    16'd4502: out <= 16'hFCAA;    16'd4503: out <= 16'h0100;
    16'd4504: out <= 16'h001B;    16'd4505: out <= 16'h027D;    16'd4506: out <= 16'h06A8;    16'd4507: out <= 16'hF7BC;
    16'd4508: out <= 16'h065C;    16'd4509: out <= 16'hFEC1;    16'd4510: out <= 16'hFF78;    16'd4511: out <= 16'hF9DD;
    16'd4512: out <= 16'hFE41;    16'd4513: out <= 16'h0517;    16'd4514: out <= 16'h09FD;    16'd4515: out <= 16'h01D2;
    16'd4516: out <= 16'hFCD9;    16'd4517: out <= 16'h093F;    16'd4518: out <= 16'hFD5B;    16'd4519: out <= 16'h047E;
    16'd4520: out <= 16'h03FE;    16'd4521: out <= 16'hFECE;    16'd4522: out <= 16'h065B;    16'd4523: out <= 16'hFDE0;
    16'd4524: out <= 16'h02EE;    16'd4525: out <= 16'h062E;    16'd4526: out <= 16'h07C5;    16'd4527: out <= 16'hFDDD;
    16'd4528: out <= 16'hFE98;    16'd4529: out <= 16'h038C;    16'd4530: out <= 16'h09A0;    16'd4531: out <= 16'h036F;
    16'd4532: out <= 16'hF9E9;    16'd4533: out <= 16'hF8AB;    16'd4534: out <= 16'hFFA5;    16'd4535: out <= 16'hFA8F;
    16'd4536: out <= 16'h0048;    16'd4537: out <= 16'hFF25;    16'd4538: out <= 16'h0290;    16'd4539: out <= 16'h03AC;
    16'd4540: out <= 16'h0394;    16'd4541: out <= 16'hFBCF;    16'd4542: out <= 16'h0311;    16'd4543: out <= 16'h00AE;
    16'd4544: out <= 16'h0099;    16'd4545: out <= 16'h0625;    16'd4546: out <= 16'hFB77;    16'd4547: out <= 16'h01EA;
    16'd4548: out <= 16'hFEF7;    16'd4549: out <= 16'h04B8;    16'd4550: out <= 16'h01EA;    16'd4551: out <= 16'h0492;
    16'd4552: out <= 16'hFAB1;    16'd4553: out <= 16'h0144;    16'd4554: out <= 16'hFFF6;    16'd4555: out <= 16'h0572;
    16'd4556: out <= 16'hFC41;    16'd4557: out <= 16'hFEC1;    16'd4558: out <= 16'h010A;    16'd4559: out <= 16'hF98F;
    16'd4560: out <= 16'hFD6C;    16'd4561: out <= 16'h0271;    16'd4562: out <= 16'h02E5;    16'd4563: out <= 16'hFD0F;
    16'd4564: out <= 16'hFC02;    16'd4565: out <= 16'h0958;    16'd4566: out <= 16'h005D;    16'd4567: out <= 16'hFE7D;
    16'd4568: out <= 16'hFD50;    16'd4569: out <= 16'hFE3F;    16'd4570: out <= 16'hFF4C;    16'd4571: out <= 16'h02AA;
    16'd4572: out <= 16'hF882;    16'd4573: out <= 16'h001A;    16'd4574: out <= 16'h0367;    16'd4575: out <= 16'h0694;
    16'd4576: out <= 16'hFED1;    16'd4577: out <= 16'hFF8E;    16'd4578: out <= 16'h06A1;    16'd4579: out <= 16'h013A;
    16'd4580: out <= 16'hFFEF;    16'd4581: out <= 16'hFD69;    16'd4582: out <= 16'hFB50;    16'd4583: out <= 16'h005A;
    16'd4584: out <= 16'hF7FD;    16'd4585: out <= 16'h06D9;    16'd4586: out <= 16'hFCBE;    16'd4587: out <= 16'h05BC;
    16'd4588: out <= 16'h0669;    16'd4589: out <= 16'hFBDE;    16'd4590: out <= 16'h00E9;    16'd4591: out <= 16'h060D;
    16'd4592: out <= 16'h0B1E;    16'd4593: out <= 16'hFB3D;    16'd4594: out <= 16'hFE43;    16'd4595: out <= 16'hFEFA;
    16'd4596: out <= 16'hFF2D;    16'd4597: out <= 16'h03E5;    16'd4598: out <= 16'hFCE6;    16'd4599: out <= 16'hFF6F;
    16'd4600: out <= 16'h0203;    16'd4601: out <= 16'h0666;    16'd4602: out <= 16'hFEAB;    16'd4603: out <= 16'hFD4C;
    16'd4604: out <= 16'hFD65;    16'd4605: out <= 16'h01EF;    16'd4606: out <= 16'h00A0;    16'd4607: out <= 16'hFE22;
    16'd4608: out <= 16'hFE8F;    16'd4609: out <= 16'hFD9D;    16'd4610: out <= 16'hF7F3;    16'd4611: out <= 16'hFB3C;
    16'd4612: out <= 16'h0100;    16'd4613: out <= 16'hFDCE;    16'd4614: out <= 16'hFAAA;    16'd4615: out <= 16'hFDEE;
    16'd4616: out <= 16'h05D4;    16'd4617: out <= 16'h0284;    16'd4618: out <= 16'h0293;    16'd4619: out <= 16'hFC25;
    16'd4620: out <= 16'h0073;    16'd4621: out <= 16'h028C;    16'd4622: out <= 16'h0152;    16'd4623: out <= 16'h0247;
    16'd4624: out <= 16'hFF13;    16'd4625: out <= 16'hF698;    16'd4626: out <= 16'h05BB;    16'd4627: out <= 16'h04C4;
    16'd4628: out <= 16'hFE1C;    16'd4629: out <= 16'h0046;    16'd4630: out <= 16'h0543;    16'd4631: out <= 16'hFCD8;
    16'd4632: out <= 16'hFA6E;    16'd4633: out <= 16'h0358;    16'd4634: out <= 16'h069D;    16'd4635: out <= 16'hFFF1;
    16'd4636: out <= 16'hFBE4;    16'd4637: out <= 16'h0109;    16'd4638: out <= 16'hFA3F;    16'd4639: out <= 16'hFB30;
    16'd4640: out <= 16'hFA98;    16'd4641: out <= 16'hFEE0;    16'd4642: out <= 16'h05F9;    16'd4643: out <= 16'h07D9;
    16'd4644: out <= 16'hFE2A;    16'd4645: out <= 16'hFDEA;    16'd4646: out <= 16'hFA29;    16'd4647: out <= 16'hFA58;
    16'd4648: out <= 16'hFB0A;    16'd4649: out <= 16'h02AB;    16'd4650: out <= 16'h08D1;    16'd4651: out <= 16'h0263;
    16'd4652: out <= 16'h039A;    16'd4653: out <= 16'h0118;    16'd4654: out <= 16'hFE1E;    16'd4655: out <= 16'hFCAA;
    16'd4656: out <= 16'h0071;    16'd4657: out <= 16'hFB19;    16'd4658: out <= 16'hFD83;    16'd4659: out <= 16'hFB32;
    16'd4660: out <= 16'h016C;    16'd4661: out <= 16'hFA8C;    16'd4662: out <= 16'hFA7D;    16'd4663: out <= 16'hF72E;
    16'd4664: out <= 16'h026D;    16'd4665: out <= 16'hFF69;    16'd4666: out <= 16'h06EB;    16'd4667: out <= 16'h0B11;
    16'd4668: out <= 16'h01A8;    16'd4669: out <= 16'h03D1;    16'd4670: out <= 16'h02D7;    16'd4671: out <= 16'h0553;
    16'd4672: out <= 16'h092A;    16'd4673: out <= 16'h0577;    16'd4674: out <= 16'h02BB;    16'd4675: out <= 16'h06C4;
    16'd4676: out <= 16'hFF3E;    16'd4677: out <= 16'h0739;    16'd4678: out <= 16'h03E3;    16'd4679: out <= 16'h053C;
    16'd4680: out <= 16'hFFDB;    16'd4681: out <= 16'h030B;    16'd4682: out <= 16'h0911;    16'd4683: out <= 16'h012C;
    16'd4684: out <= 16'h028C;    16'd4685: out <= 16'h0B43;    16'd4686: out <= 16'h017E;    16'd4687: out <= 16'h0179;
    16'd4688: out <= 16'h0658;    16'd4689: out <= 16'hFC22;    16'd4690: out <= 16'h0273;    16'd4691: out <= 16'h0A6C;
    16'd4692: out <= 16'h04CC;    16'd4693: out <= 16'h0352;    16'd4694: out <= 16'h053B;    16'd4695: out <= 16'h051E;
    16'd4696: out <= 16'hFFC4;    16'd4697: out <= 16'h02B4;    16'd4698: out <= 16'hFFCB;    16'd4699: out <= 16'h0A3C;
    16'd4700: out <= 16'h08DE;    16'd4701: out <= 16'h00BB;    16'd4702: out <= 16'hFDCF;    16'd4703: out <= 16'h01D5;
    16'd4704: out <= 16'h07AB;    16'd4705: out <= 16'h046F;    16'd4706: out <= 16'h0264;    16'd4707: out <= 16'h0090;
    16'd4708: out <= 16'hFEB7;    16'd4709: out <= 16'h07CD;    16'd4710: out <= 16'h0523;    16'd4711: out <= 16'h0571;
    16'd4712: out <= 16'h052A;    16'd4713: out <= 16'hFFA5;    16'd4714: out <= 16'h02B8;    16'd4715: out <= 16'h0386;
    16'd4716: out <= 16'h010B;    16'd4717: out <= 16'h0E14;    16'd4718: out <= 16'h03B0;    16'd4719: out <= 16'h04D6;
    16'd4720: out <= 16'h04F3;    16'd4721: out <= 16'h0A4B;    16'd4722: out <= 16'h02E3;    16'd4723: out <= 16'h0CF4;
    16'd4724: out <= 16'h0278;    16'd4725: out <= 16'h0094;    16'd4726: out <= 16'h0504;    16'd4727: out <= 16'h0040;
    16'd4728: out <= 16'h02A0;    16'd4729: out <= 16'h029A;    16'd4730: out <= 16'h02F2;    16'd4731: out <= 16'h09C1;
    16'd4732: out <= 16'h07FD;    16'd4733: out <= 16'h0718;    16'd4734: out <= 16'hFB2D;    16'd4735: out <= 16'h0819;
    16'd4736: out <= 16'h06B0;    16'd4737: out <= 16'h037F;    16'd4738: out <= 16'hFF0B;    16'd4739: out <= 16'h05E1;
    16'd4740: out <= 16'h0643;    16'd4741: out <= 16'h01C8;    16'd4742: out <= 16'h081F;    16'd4743: out <= 16'h01F2;
    16'd4744: out <= 16'h0222;    16'd4745: out <= 16'h00DC;    16'd4746: out <= 16'h0143;    16'd4747: out <= 16'h04AB;
    16'd4748: out <= 16'h02F8;    16'd4749: out <= 16'h05C6;    16'd4750: out <= 16'h056F;    16'd4751: out <= 16'h028E;
    16'd4752: out <= 16'h06FB;    16'd4753: out <= 16'h0619;    16'd4754: out <= 16'h05F7;    16'd4755: out <= 16'h06E7;
    16'd4756: out <= 16'h02FF;    16'd4757: out <= 16'h03ED;    16'd4758: out <= 16'h007A;    16'd4759: out <= 16'h0153;
    16'd4760: out <= 16'hFC3E;    16'd4761: out <= 16'h0794;    16'd4762: out <= 16'h05F3;    16'd4763: out <= 16'h0919;
    16'd4764: out <= 16'h03C9;    16'd4765: out <= 16'h09E7;    16'd4766: out <= 16'hFB76;    16'd4767: out <= 16'h0929;
    16'd4768: out <= 16'h051C;    16'd4769: out <= 16'h022F;    16'd4770: out <= 16'h06EA;    16'd4771: out <= 16'h05F1;
    16'd4772: out <= 16'h0381;    16'd4773: out <= 16'h026A;    16'd4774: out <= 16'h09AA;    16'd4775: out <= 16'h090F;
    16'd4776: out <= 16'h0AA0;    16'd4777: out <= 16'hFE76;    16'd4778: out <= 16'h0020;    16'd4779: out <= 16'h0554;
    16'd4780: out <= 16'h0259;    16'd4781: out <= 16'h098E;    16'd4782: out <= 16'h05D9;    16'd4783: out <= 16'h0E13;
    16'd4784: out <= 16'h008E;    16'd4785: out <= 16'h07D1;    16'd4786: out <= 16'hFFFB;    16'd4787: out <= 16'h090E;
    16'd4788: out <= 16'h0362;    16'd4789: out <= 16'h07A0;    16'd4790: out <= 16'h0721;    16'd4791: out <= 16'h051A;
    16'd4792: out <= 16'h0440;    16'd4793: out <= 16'h02BA;    16'd4794: out <= 16'h02B5;    16'd4795: out <= 16'hFDF3;
    16'd4796: out <= 16'hF89D;    16'd4797: out <= 16'hFAEF;    16'd4798: out <= 16'h041F;    16'd4799: out <= 16'hFB08;
    16'd4800: out <= 16'hFDB5;    16'd4801: out <= 16'h0590;    16'd4802: out <= 16'h0080;    16'd4803: out <= 16'hFCAB;
    16'd4804: out <= 16'h01A7;    16'd4805: out <= 16'hFCCD;    16'd4806: out <= 16'h0127;    16'd4807: out <= 16'hFC68;
    16'd4808: out <= 16'hFD55;    16'd4809: out <= 16'h02C4;    16'd4810: out <= 16'hF893;    16'd4811: out <= 16'hFCE2;
    16'd4812: out <= 16'h00EC;    16'd4813: out <= 16'h0388;    16'd4814: out <= 16'h02DF;    16'd4815: out <= 16'hFCDD;
    16'd4816: out <= 16'hFF86;    16'd4817: out <= 16'hFBE0;    16'd4818: out <= 16'h049B;    16'd4819: out <= 16'hFD69;
    16'd4820: out <= 16'hFF8A;    16'd4821: out <= 16'h011A;    16'd4822: out <= 16'h0388;    16'd4823: out <= 16'h0302;
    16'd4824: out <= 16'hFCAD;    16'd4825: out <= 16'h0115;    16'd4826: out <= 16'hFB9A;    16'd4827: out <= 16'hFD2E;
    16'd4828: out <= 16'h046B;    16'd4829: out <= 16'hFF36;    16'd4830: out <= 16'h051D;    16'd4831: out <= 16'h01FB;
    16'd4832: out <= 16'h0382;    16'd4833: out <= 16'hFEB6;    16'd4834: out <= 16'h01A4;    16'd4835: out <= 16'h03BA;
    16'd4836: out <= 16'hFF56;    16'd4837: out <= 16'h026E;    16'd4838: out <= 16'hFD2C;    16'd4839: out <= 16'h00B6;
    16'd4840: out <= 16'hFF32;    16'd4841: out <= 16'h02AB;    16'd4842: out <= 16'hFBF2;    16'd4843: out <= 16'h0576;
    16'd4844: out <= 16'h0252;    16'd4845: out <= 16'h071F;    16'd4846: out <= 16'hF724;    16'd4847: out <= 16'hFC6C;
    16'd4848: out <= 16'h0387;    16'd4849: out <= 16'h0431;    16'd4850: out <= 16'h029C;    16'd4851: out <= 16'h03A6;
    16'd4852: out <= 16'hFE6B;    16'd4853: out <= 16'h0104;    16'd4854: out <= 16'hFC15;    16'd4855: out <= 16'h0100;
    16'd4856: out <= 16'h0255;    16'd4857: out <= 16'h038A;    16'd4858: out <= 16'h03B5;    16'd4859: out <= 16'hFF9E;
    16'd4860: out <= 16'hF5CA;    16'd4861: out <= 16'h045E;    16'd4862: out <= 16'hFC85;    16'd4863: out <= 16'h00A6;
    16'd4864: out <= 16'h00B0;    16'd4865: out <= 16'hFFA5;    16'd4866: out <= 16'hFA2C;    16'd4867: out <= 16'h065F;
    16'd4868: out <= 16'hFD2B;    16'd4869: out <= 16'h01B0;    16'd4870: out <= 16'h0263;    16'd4871: out <= 16'h010A;
    16'd4872: out <= 16'h0030;    16'd4873: out <= 16'h0247;    16'd4874: out <= 16'h006C;    16'd4875: out <= 16'hFF51;
    16'd4876: out <= 16'h0464;    16'd4877: out <= 16'h08A2;    16'd4878: out <= 16'h08DF;    16'd4879: out <= 16'hF7E1;
    16'd4880: out <= 16'hFDCD;    16'd4881: out <= 16'h071F;    16'd4882: out <= 16'hFD7C;    16'd4883: out <= 16'h020B;
    16'd4884: out <= 16'hFE39;    16'd4885: out <= 16'hF9FE;    16'd4886: out <= 16'h009C;    16'd4887: out <= 16'h0194;
    16'd4888: out <= 16'h029D;    16'd4889: out <= 16'h0149;    16'd4890: out <= 16'hFC57;    16'd4891: out <= 16'hFEFF;
    16'd4892: out <= 16'h0297;    16'd4893: out <= 16'h04E2;    16'd4894: out <= 16'h068D;    16'd4895: out <= 16'hFF3C;
    16'd4896: out <= 16'h0165;    16'd4897: out <= 16'hFEAC;    16'd4898: out <= 16'hFA83;    16'd4899: out <= 16'h047A;
    16'd4900: out <= 16'h03A1;    16'd4901: out <= 16'hFF85;    16'd4902: out <= 16'hFB9B;    16'd4903: out <= 16'hFC75;
    16'd4904: out <= 16'hFC2D;    16'd4905: out <= 16'h045F;    16'd4906: out <= 16'hFF79;    16'd4907: out <= 16'h01DE;
    16'd4908: out <= 16'h04F0;    16'd4909: out <= 16'hF650;    16'd4910: out <= 16'hFD3F;    16'd4911: out <= 16'h033D;
    16'd4912: out <= 16'h03A0;    16'd4913: out <= 16'hFDB2;    16'd4914: out <= 16'hFA39;    16'd4915: out <= 16'hFDFF;
    16'd4916: out <= 16'h01CA;    16'd4917: out <= 16'h0604;    16'd4918: out <= 16'hFF9C;    16'd4919: out <= 16'h0897;
    16'd4920: out <= 16'hFCD6;    16'd4921: out <= 16'h02C8;    16'd4922: out <= 16'h07E8;    16'd4923: out <= 16'h038D;
    16'd4924: out <= 16'h02BB;    16'd4925: out <= 16'h055B;    16'd4926: out <= 16'h0B5E;    16'd4927: out <= 16'h09DF;
    16'd4928: out <= 16'hFDA3;    16'd4929: out <= 16'h0021;    16'd4930: out <= 16'h046C;    16'd4931: out <= 16'h033B;
    16'd4932: out <= 16'h033A;    16'd4933: out <= 16'h088E;    16'd4934: out <= 16'h02AB;    16'd4935: out <= 16'h0716;
    16'd4936: out <= 16'h060C;    16'd4937: out <= 16'h0BD2;    16'd4938: out <= 16'h03C4;    16'd4939: out <= 16'h070A;
    16'd4940: out <= 16'h097D;    16'd4941: out <= 16'hFE7D;    16'd4942: out <= 16'h024D;    16'd4943: out <= 16'h082B;
    16'd4944: out <= 16'h0AE1;    16'd4945: out <= 16'hFEA6;    16'd4946: out <= 16'h0487;    16'd4947: out <= 16'h0558;
    16'd4948: out <= 16'h0445;    16'd4949: out <= 16'h0361;    16'd4950: out <= 16'h0666;    16'd4951: out <= 16'h0855;
    16'd4952: out <= 16'h01D9;    16'd4953: out <= 16'h0365;    16'd4954: out <= 16'h0948;    16'd4955: out <= 16'h06D9;
    16'd4956: out <= 16'h0253;    16'd4957: out <= 16'h033A;    16'd4958: out <= 16'hFB75;    16'd4959: out <= 16'h0B3D;
    16'd4960: out <= 16'h03A4;    16'd4961: out <= 16'hFF79;    16'd4962: out <= 16'h03E8;    16'd4963: out <= 16'hFD1A;
    16'd4964: out <= 16'h0716;    16'd4965: out <= 16'h03A1;    16'd4966: out <= 16'hFDDB;    16'd4967: out <= 16'h01F1;
    16'd4968: out <= 16'hFE84;    16'd4969: out <= 16'h01BF;    16'd4970: out <= 16'h03BC;    16'd4971: out <= 16'h0272;
    16'd4972: out <= 16'h05C4;    16'd4973: out <= 16'h057E;    16'd4974: out <= 16'h0336;    16'd4975: out <= 16'h0566;
    16'd4976: out <= 16'hFFE9;    16'd4977: out <= 16'h08E1;    16'd4978: out <= 16'h0235;    16'd4979: out <= 16'hFAF9;
    16'd4980: out <= 16'hFEE6;    16'd4981: out <= 16'h0BE9;    16'd4982: out <= 16'h04EF;    16'd4983: out <= 16'h0794;
    16'd4984: out <= 16'h08A6;    16'd4985: out <= 16'h0457;    16'd4986: out <= 16'hFF11;    16'd4987: out <= 16'h0086;
    16'd4988: out <= 16'h01F1;    16'd4989: out <= 16'h06CE;    16'd4990: out <= 16'h0905;    16'd4991: out <= 16'hFB64;
    16'd4992: out <= 16'h0108;    16'd4993: out <= 16'h0940;    16'd4994: out <= 16'h0AC8;    16'd4995: out <= 16'h0473;
    16'd4996: out <= 16'h0800;    16'd4997: out <= 16'h0154;    16'd4998: out <= 16'hFEEC;    16'd4999: out <= 16'h0223;
    16'd5000: out <= 16'hFF14;    16'd5001: out <= 16'h0941;    16'd5002: out <= 16'h0399;    16'd5003: out <= 16'hFE80;
    16'd5004: out <= 16'h0418;    16'd5005: out <= 16'h06B0;    16'd5006: out <= 16'h0BA1;    16'd5007: out <= 16'h0559;
    16'd5008: out <= 16'h0762;    16'd5009: out <= 16'h0221;    16'd5010: out <= 16'h0348;    16'd5011: out <= 16'h019A;
    16'd5012: out <= 16'h0697;    16'd5013: out <= 16'h0E0E;    16'd5014: out <= 16'h0072;    16'd5015: out <= 16'h06F6;
    16'd5016: out <= 16'h03BF;    16'd5017: out <= 16'h06D8;    16'd5018: out <= 16'h04F4;    16'd5019: out <= 16'h0DA0;
    16'd5020: out <= 16'hFECB;    16'd5021: out <= 16'hFF23;    16'd5022: out <= 16'h0426;    16'd5023: out <= 16'h04EE;
    16'd5024: out <= 16'hFFA8;    16'd5025: out <= 16'h03DE;    16'd5026: out <= 16'h07EF;    16'd5027: out <= 16'h030A;
    16'd5028: out <= 16'hFD69;    16'd5029: out <= 16'h00D1;    16'd5030: out <= 16'h01CE;    16'd5031: out <= 16'hFEB0;
    16'd5032: out <= 16'h0A46;    16'd5033: out <= 16'h05A8;    16'd5034: out <= 16'h0250;    16'd5035: out <= 16'h0186;
    16'd5036: out <= 16'hFD84;    16'd5037: out <= 16'hFCA4;    16'd5038: out <= 16'h049C;    16'd5039: out <= 16'h0345;
    16'd5040: out <= 16'hFDA4;    16'd5041: out <= 16'h0B9D;    16'd5042: out <= 16'h02E8;    16'd5043: out <= 16'h05FA;
    16'd5044: out <= 16'h074D;    16'd5045: out <= 16'h0E33;    16'd5046: out <= 16'h0861;    16'd5047: out <= 16'h0169;
    16'd5048: out <= 16'h017C;    16'd5049: out <= 16'h0707;    16'd5050: out <= 16'hFEC3;    16'd5051: out <= 16'h0097;
    16'd5052: out <= 16'hFACF;    16'd5053: out <= 16'h03AF;    16'd5054: out <= 16'h009C;    16'd5055: out <= 16'h043B;
    16'd5056: out <= 16'hFC80;    16'd5057: out <= 16'h038C;    16'd5058: out <= 16'h073E;    16'd5059: out <= 16'hFB48;
    16'd5060: out <= 16'hFAE0;    16'd5061: out <= 16'h04D4;    16'd5062: out <= 16'h0439;    16'd5063: out <= 16'h013D;
    16'd5064: out <= 16'h00DA;    16'd5065: out <= 16'h02A9;    16'd5066: out <= 16'h013B;    16'd5067: out <= 16'hFC7A;
    16'd5068: out <= 16'hFA2E;    16'd5069: out <= 16'hFF18;    16'd5070: out <= 16'h0299;    16'd5071: out <= 16'hFE2E;
    16'd5072: out <= 16'h0895;    16'd5073: out <= 16'h043F;    16'd5074: out <= 16'h00FB;    16'd5075: out <= 16'h027A;
    16'd5076: out <= 16'hFFBD;    16'd5077: out <= 16'h0023;    16'd5078: out <= 16'h02F0;    16'd5079: out <= 16'h0031;
    16'd5080: out <= 16'h0483;    16'd5081: out <= 16'hFCC0;    16'd5082: out <= 16'hF97D;    16'd5083: out <= 16'h0277;
    16'd5084: out <= 16'h012A;    16'd5085: out <= 16'h0518;    16'd5086: out <= 16'hFEAC;    16'd5087: out <= 16'hFA23;
    16'd5088: out <= 16'h07F2;    16'd5089: out <= 16'hFD38;    16'd5090: out <= 16'h03BB;    16'd5091: out <= 16'h00F4;
    16'd5092: out <= 16'h003A;    16'd5093: out <= 16'h0304;    16'd5094: out <= 16'h0355;    16'd5095: out <= 16'h0221;
    16'd5096: out <= 16'hFD89;    16'd5097: out <= 16'h007D;    16'd5098: out <= 16'h0112;    16'd5099: out <= 16'h0020;
    16'd5100: out <= 16'h040D;    16'd5101: out <= 16'hFCA2;    16'd5102: out <= 16'h094A;    16'd5103: out <= 16'h071E;
    16'd5104: out <= 16'hFE1B;    16'd5105: out <= 16'h0458;    16'd5106: out <= 16'h040E;    16'd5107: out <= 16'h051C;
    16'd5108: out <= 16'hF7B5;    16'd5109: out <= 16'h012C;    16'd5110: out <= 16'hFF89;    16'd5111: out <= 16'h00E4;
    16'd5112: out <= 16'h0609;    16'd5113: out <= 16'hFDC6;    16'd5114: out <= 16'hFAB8;    16'd5115: out <= 16'hFED6;
    16'd5116: out <= 16'hFBDA;    16'd5117: out <= 16'h02CC;    16'd5118: out <= 16'h00CC;    16'd5119: out <= 16'h00F4;
    16'd5120: out <= 16'hF852;    16'd5121: out <= 16'hFABE;    16'd5122: out <= 16'hFB67;    16'd5123: out <= 16'hFF4D;
    16'd5124: out <= 16'h0352;    16'd5125: out <= 16'h02B5;    16'd5126: out <= 16'h02D0;    16'd5127: out <= 16'hF838;
    16'd5128: out <= 16'h046A;    16'd5129: out <= 16'hFED5;    16'd5130: out <= 16'hFC37;    16'd5131: out <= 16'h008C;
    16'd5132: out <= 16'h0015;    16'd5133: out <= 16'h0049;    16'd5134: out <= 16'hFB58;    16'd5135: out <= 16'hFC99;
    16'd5136: out <= 16'h00B9;    16'd5137: out <= 16'h02F9;    16'd5138: out <= 16'h006D;    16'd5139: out <= 16'hFE22;
    16'd5140: out <= 16'hFFBF;    16'd5141: out <= 16'hFE94;    16'd5142: out <= 16'hFB06;    16'd5143: out <= 16'h02A2;
    16'd5144: out <= 16'h038C;    16'd5145: out <= 16'h02A9;    16'd5146: out <= 16'hFE99;    16'd5147: out <= 16'hFD43;
    16'd5148: out <= 16'hFD54;    16'd5149: out <= 16'hFC91;    16'd5150: out <= 16'h0124;    16'd5151: out <= 16'hFFB6;
    16'd5152: out <= 16'h04CA;    16'd5153: out <= 16'hFE54;    16'd5154: out <= 16'hFE3B;    16'd5155: out <= 16'h0096;
    16'd5156: out <= 16'hFEA8;    16'd5157: out <= 16'hFF39;    16'd5158: out <= 16'hFF68;    16'd5159: out <= 16'h006F;
    16'd5160: out <= 16'hFF0D;    16'd5161: out <= 16'hF5A1;    16'd5162: out <= 16'hFDEC;    16'd5163: out <= 16'hFFFB;
    16'd5164: out <= 16'hFEBD;    16'd5165: out <= 16'hFAF3;    16'd5166: out <= 16'h0277;    16'd5167: out <= 16'h0050;
    16'd5168: out <= 16'hFB6C;    16'd5169: out <= 16'h00CA;    16'd5170: out <= 16'hFE7D;    16'd5171: out <= 16'hFDE6;
    16'd5172: out <= 16'hFFBD;    16'd5173: out <= 16'h0180;    16'd5174: out <= 16'hFC5E;    16'd5175: out <= 16'h05F3;
    16'd5176: out <= 16'h02CA;    16'd5177: out <= 16'hFEE4;    16'd5178: out <= 16'h0631;    16'd5179: out <= 16'h00E8;
    16'd5180: out <= 16'h04D3;    16'd5181: out <= 16'hFD86;    16'd5182: out <= 16'h045B;    16'd5183: out <= 16'hFDD9;
    16'd5184: out <= 16'h0924;    16'd5185: out <= 16'hFEB0;    16'd5186: out <= 16'h0628;    16'd5187: out <= 16'h077F;
    16'd5188: out <= 16'h0496;    16'd5189: out <= 16'h04B8;    16'd5190: out <= 16'h0B78;    16'd5191: out <= 16'h0472;
    16'd5192: out <= 16'h0897;    16'd5193: out <= 16'hFBA2;    16'd5194: out <= 16'h0C6A;    16'd5195: out <= 16'h07B2;
    16'd5196: out <= 16'h06D7;    16'd5197: out <= 16'h087F;    16'd5198: out <= 16'h080D;    16'd5199: out <= 16'h031E;
    16'd5200: out <= 16'h04A3;    16'd5201: out <= 16'h011F;    16'd5202: out <= 16'h02A7;    16'd5203: out <= 16'h0A0E;
    16'd5204: out <= 16'h0355;    16'd5205: out <= 16'h0920;    16'd5206: out <= 16'h0069;    16'd5207: out <= 16'h028B;
    16'd5208: out <= 16'h02DE;    16'd5209: out <= 16'h00CD;    16'd5210: out <= 16'h0906;    16'd5211: out <= 16'h0E85;
    16'd5212: out <= 16'h05E9;    16'd5213: out <= 16'h03C4;    16'd5214: out <= 16'h0790;    16'd5215: out <= 16'h097B;
    16'd5216: out <= 16'h0530;    16'd5217: out <= 16'h0823;    16'd5218: out <= 16'h0199;    16'd5219: out <= 16'h05EF;
    16'd5220: out <= 16'h04AF;    16'd5221: out <= 16'h0380;    16'd5222: out <= 16'h09F4;    16'd5223: out <= 16'h079C;
    16'd5224: out <= 16'h04F8;    16'd5225: out <= 16'h078F;    16'd5226: out <= 16'hFBAD;    16'd5227: out <= 16'h030C;
    16'd5228: out <= 16'h0459;    16'd5229: out <= 16'h0981;    16'd5230: out <= 16'h05BB;    16'd5231: out <= 16'h04B2;
    16'd5232: out <= 16'h0429;    16'd5233: out <= 16'h033C;    16'd5234: out <= 16'hFEB9;    16'd5235: out <= 16'h025E;
    16'd5236: out <= 16'hFBF5;    16'd5237: out <= 16'h04AC;    16'd5238: out <= 16'h0240;    16'd5239: out <= 16'h032D;
    16'd5240: out <= 16'h0307;    16'd5241: out <= 16'h048E;    16'd5242: out <= 16'h0056;    16'd5243: out <= 16'hFFED;
    16'd5244: out <= 16'h04AB;    16'd5245: out <= 16'h03B4;    16'd5246: out <= 16'h06A4;    16'd5247: out <= 16'h095A;
    16'd5248: out <= 16'h02C7;    16'd5249: out <= 16'h0415;    16'd5250: out <= 16'h051A;    16'd5251: out <= 16'h039E;
    16'd5252: out <= 16'h0024;    16'd5253: out <= 16'hFE7E;    16'd5254: out <= 16'h048E;    16'd5255: out <= 16'h065F;
    16'd5256: out <= 16'h06FD;    16'd5257: out <= 16'h0D5F;    16'd5258: out <= 16'h0943;    16'd5259: out <= 16'hFEAF;
    16'd5260: out <= 16'h02D3;    16'd5261: out <= 16'h061D;    16'd5262: out <= 16'h0995;    16'd5263: out <= 16'h00BB;
    16'd5264: out <= 16'h0945;    16'd5265: out <= 16'h06E1;    16'd5266: out <= 16'h0230;    16'd5267: out <= 16'hFE55;
    16'd5268: out <= 16'h0027;    16'd5269: out <= 16'h0127;    16'd5270: out <= 16'h04CD;    16'd5271: out <= 16'h022F;
    16'd5272: out <= 16'h03CC;    16'd5273: out <= 16'h0338;    16'd5274: out <= 16'h0542;    16'd5275: out <= 16'h0844;
    16'd5276: out <= 16'h0B66;    16'd5277: out <= 16'h0C90;    16'd5278: out <= 16'h030E;    16'd5279: out <= 16'h0876;
    16'd5280: out <= 16'h036A;    16'd5281: out <= 16'h0328;    16'd5282: out <= 16'hFCD9;    16'd5283: out <= 16'h0CDB;
    16'd5284: out <= 16'h0331;    16'd5285: out <= 16'h02B5;    16'd5286: out <= 16'h0711;    16'd5287: out <= 16'hFFFD;
    16'd5288: out <= 16'h02E4;    16'd5289: out <= 16'h0783;    16'd5290: out <= 16'hFA35;    16'd5291: out <= 16'h0165;
    16'd5292: out <= 16'h0111;    16'd5293: out <= 16'h0454;    16'd5294: out <= 16'h0200;    16'd5295: out <= 16'h06A8;
    16'd5296: out <= 16'h00C3;    16'd5297: out <= 16'h0512;    16'd5298: out <= 16'h0148;    16'd5299: out <= 16'hFE0F;
    16'd5300: out <= 16'h0DA4;    16'd5301: out <= 16'h07CB;    16'd5302: out <= 16'hFFF2;    16'd5303: out <= 16'h03AA;
    16'd5304: out <= 16'hFC4C;    16'd5305: out <= 16'h0058;    16'd5306: out <= 16'h0228;    16'd5307: out <= 16'h074C;
    16'd5308: out <= 16'h01CB;    16'd5309: out <= 16'hFCC1;    16'd5310: out <= 16'hFFC1;    16'd5311: out <= 16'hFC7D;
    16'd5312: out <= 16'hFEB4;    16'd5313: out <= 16'h04B3;    16'd5314: out <= 16'hFED1;    16'd5315: out <= 16'hF8AD;
    16'd5316: out <= 16'h01F6;    16'd5317: out <= 16'h014F;    16'd5318: out <= 16'h016B;    16'd5319: out <= 16'h0644;
    16'd5320: out <= 16'hFFA8;    16'd5321: out <= 16'hFF06;    16'd5322: out <= 16'h037E;    16'd5323: out <= 16'hFCF8;
    16'd5324: out <= 16'hFD45;    16'd5325: out <= 16'hFAEC;    16'd5326: out <= 16'h009E;    16'd5327: out <= 16'h0080;
    16'd5328: out <= 16'hFC05;    16'd5329: out <= 16'h05EF;    16'd5330: out <= 16'h06E3;    16'd5331: out <= 16'hFFEE;
    16'd5332: out <= 16'hFF9B;    16'd5333: out <= 16'h01A2;    16'd5334: out <= 16'h0525;    16'd5335: out <= 16'h04BF;
    16'd5336: out <= 16'h0353;    16'd5337: out <= 16'hFE4C;    16'd5338: out <= 16'hFA9D;    16'd5339: out <= 16'h04E0;
    16'd5340: out <= 16'h00FF;    16'd5341: out <= 16'h006F;    16'd5342: out <= 16'hFC11;    16'd5343: out <= 16'h022F;
    16'd5344: out <= 16'hFE1A;    16'd5345: out <= 16'hFAD3;    16'd5346: out <= 16'h0453;    16'd5347: out <= 16'h0149;
    16'd5348: out <= 16'h0150;    16'd5349: out <= 16'h03CA;    16'd5350: out <= 16'hF9E5;    16'd5351: out <= 16'h0615;
    16'd5352: out <= 16'hFDC7;    16'd5353: out <= 16'h0305;    16'd5354: out <= 16'h006B;    16'd5355: out <= 16'hFD66;
    16'd5356: out <= 16'h0096;    16'd5357: out <= 16'h0111;    16'd5358: out <= 16'h002E;    16'd5359: out <= 16'h0368;
    16'd5360: out <= 16'h0178;    16'd5361: out <= 16'h0078;    16'd5362: out <= 16'hF90E;    16'd5363: out <= 16'h00EB;
    16'd5364: out <= 16'h0516;    16'd5365: out <= 16'hFCBC;    16'd5366: out <= 16'h05B1;    16'd5367: out <= 16'hFFA9;
    16'd5368: out <= 16'hFF6F;    16'd5369: out <= 16'hFD00;    16'd5370: out <= 16'hF902;    16'd5371: out <= 16'h0733;
    16'd5372: out <= 16'h027E;    16'd5373: out <= 16'h0382;    16'd5374: out <= 16'hFFF8;    16'd5375: out <= 16'hFC10;
    16'd5376: out <= 16'h0047;    16'd5377: out <= 16'h0536;    16'd5378: out <= 16'hFC2F;    16'd5379: out <= 16'hFC33;
    16'd5380: out <= 16'hFE1D;    16'd5381: out <= 16'hFCC4;    16'd5382: out <= 16'hFBE8;    16'd5383: out <= 16'hFE71;
    16'd5384: out <= 16'h01F8;    16'd5385: out <= 16'hFEB4;    16'd5386: out <= 16'hFCF1;    16'd5387: out <= 16'h0176;
    16'd5388: out <= 16'hFEE0;    16'd5389: out <= 16'h0066;    16'd5390: out <= 16'hFBEF;    16'd5391: out <= 16'hFC75;
    16'd5392: out <= 16'hF9D9;    16'd5393: out <= 16'hFDE0;    16'd5394: out <= 16'h0087;    16'd5395: out <= 16'hF9C7;
    16'd5396: out <= 16'hFF3F;    16'd5397: out <= 16'h02B7;    16'd5398: out <= 16'hF864;    16'd5399: out <= 16'h0584;
    16'd5400: out <= 16'h003F;    16'd5401: out <= 16'hF838;    16'd5402: out <= 16'hFCCE;    16'd5403: out <= 16'h02BB;
    16'd5404: out <= 16'h0165;    16'd5405: out <= 16'h0054;    16'd5406: out <= 16'h01C6;    16'd5407: out <= 16'hFF09;
    16'd5408: out <= 16'hF7CC;    16'd5409: out <= 16'hFDB9;    16'd5410: out <= 16'h052B;    16'd5411: out <= 16'hFEC5;
    16'd5412: out <= 16'h05A2;    16'd5413: out <= 16'h04B7;    16'd5414: out <= 16'hFFD4;    16'd5415: out <= 16'h0412;
    16'd5416: out <= 16'hFFCC;    16'd5417: out <= 16'h048D;    16'd5418: out <= 16'hFC2F;    16'd5419: out <= 16'hFFD4;
    16'd5420: out <= 16'hFFC5;    16'd5421: out <= 16'hFD9B;    16'd5422: out <= 16'h0408;    16'd5423: out <= 16'h0300;
    16'd5424: out <= 16'h00EB;    16'd5425: out <= 16'hFF63;    16'd5426: out <= 16'hFDB6;    16'd5427: out <= 16'h04C5;
    16'd5428: out <= 16'h03AD;    16'd5429: out <= 16'h0408;    16'd5430: out <= 16'h00EF;    16'd5431: out <= 16'h0E56;
    16'd5432: out <= 16'hFF84;    16'd5433: out <= 16'hFEB0;    16'd5434: out <= 16'hFE19;    16'd5435: out <= 16'h0A13;
    16'd5436: out <= 16'h039D;    16'd5437: out <= 16'h0140;    16'd5438: out <= 16'h0283;    16'd5439: out <= 16'h020E;
    16'd5440: out <= 16'h0478;    16'd5441: out <= 16'h04EF;    16'd5442: out <= 16'h00D7;    16'd5443: out <= 16'h0754;
    16'd5444: out <= 16'h053A;    16'd5445: out <= 16'h02B4;    16'd5446: out <= 16'h0022;    16'd5447: out <= 16'h1004;
    16'd5448: out <= 16'h0396;    16'd5449: out <= 16'h0806;    16'd5450: out <= 16'h03A1;    16'd5451: out <= 16'h0406;
    16'd5452: out <= 16'h0242;    16'd5453: out <= 16'h0122;    16'd5454: out <= 16'hFE31;    16'd5455: out <= 16'h06A7;
    16'd5456: out <= 16'h0192;    16'd5457: out <= 16'h0550;    16'd5458: out <= 16'h045C;    16'd5459: out <= 16'h0654;
    16'd5460: out <= 16'h0008;    16'd5461: out <= 16'h000D;    16'd5462: out <= 16'hFA13;    16'd5463: out <= 16'h09E9;
    16'd5464: out <= 16'h0224;    16'd5465: out <= 16'h0755;    16'd5466: out <= 16'h04EB;    16'd5467: out <= 16'hFD2F;
    16'd5468: out <= 16'h03E7;    16'd5469: out <= 16'h0278;    16'd5470: out <= 16'h04A1;    16'd5471: out <= 16'h012B;
    16'd5472: out <= 16'h0634;    16'd5473: out <= 16'h0179;    16'd5474: out <= 16'h0284;    16'd5475: out <= 16'h0114;
    16'd5476: out <= 16'h069C;    16'd5477: out <= 16'h0575;    16'd5478: out <= 16'hFCA5;    16'd5479: out <= 16'h09DB;
    16'd5480: out <= 16'h0388;    16'd5481: out <= 16'hFD8C;    16'd5482: out <= 16'hFCB3;    16'd5483: out <= 16'h010D;
    16'd5484: out <= 16'h01AB;    16'd5485: out <= 16'h05A0;    16'd5486: out <= 16'h07E0;    16'd5487: out <= 16'h063D;
    16'd5488: out <= 16'h0350;    16'd5489: out <= 16'hFD3B;    16'd5490: out <= 16'h0C5C;    16'd5491: out <= 16'h03ED;
    16'd5492: out <= 16'h049B;    16'd5493: out <= 16'h0769;    16'd5494: out <= 16'h02CA;    16'd5495: out <= 16'h0514;
    16'd5496: out <= 16'h072B;    16'd5497: out <= 16'h025C;    16'd5498: out <= 16'h00AE;    16'd5499: out <= 16'hFDFA;
    16'd5500: out <= 16'h06CE;    16'd5501: out <= 16'hFE58;    16'd5502: out <= 16'h051D;    16'd5503: out <= 16'hFF55;
    16'd5504: out <= 16'h01F6;    16'd5505: out <= 16'h02D6;    16'd5506: out <= 16'h08E8;    16'd5507: out <= 16'h0640;
    16'd5508: out <= 16'h0623;    16'd5509: out <= 16'h09C9;    16'd5510: out <= 16'h05FD;    16'd5511: out <= 16'h0801;
    16'd5512: out <= 16'hFA65;    16'd5513: out <= 16'h04A0;    16'd5514: out <= 16'h03FE;    16'd5515: out <= 16'h0896;
    16'd5516: out <= 16'h014E;    16'd5517: out <= 16'h0072;    16'd5518: out <= 16'h0392;    16'd5519: out <= 16'hF9A2;
    16'd5520: out <= 16'h03EF;    16'd5521: out <= 16'h054F;    16'd5522: out <= 16'h0220;    16'd5523: out <= 16'h0273;
    16'd5524: out <= 16'h00A1;    16'd5525: out <= 16'h01FD;    16'd5526: out <= 16'h061D;    16'd5527: out <= 16'h028C;
    16'd5528: out <= 16'h0661;    16'd5529: out <= 16'h0265;    16'd5530: out <= 16'hFDE4;    16'd5531: out <= 16'h027C;
    16'd5532: out <= 16'hFFD1;    16'd5533: out <= 16'h04FC;    16'd5534: out <= 16'hFF4A;    16'd5535: out <= 16'h0100;
    16'd5536: out <= 16'h02F0;    16'd5537: out <= 16'h015A;    16'd5538: out <= 16'h0669;    16'd5539: out <= 16'h01D7;
    16'd5540: out <= 16'h094A;    16'd5541: out <= 16'hFD62;    16'd5542: out <= 16'hFF02;    16'd5543: out <= 16'h08C3;
    16'd5544: out <= 16'h062E;    16'd5545: out <= 16'h00F4;    16'd5546: out <= 16'h0801;    16'd5547: out <= 16'h011F;
    16'd5548: out <= 16'h06EE;    16'd5549: out <= 16'h02D7;    16'd5550: out <= 16'hFDF9;    16'd5551: out <= 16'h06F8;
    16'd5552: out <= 16'h082F;    16'd5553: out <= 16'hFD9F;    16'd5554: out <= 16'h012D;    16'd5555: out <= 16'h00B8;
    16'd5556: out <= 16'h00E8;    16'd5557: out <= 16'h056D;    16'd5558: out <= 16'h012A;    16'd5559: out <= 16'h0B20;
    16'd5560: out <= 16'h06FC;    16'd5561: out <= 16'h04BF;    16'd5562: out <= 16'h01DA;    16'd5563: out <= 16'h0469;
    16'd5564: out <= 16'h05D1;    16'd5565: out <= 16'hFF46;    16'd5566: out <= 16'hFED0;    16'd5567: out <= 16'hFE69;
    16'd5568: out <= 16'h03C4;    16'd5569: out <= 16'h0184;    16'd5570: out <= 16'h02C7;    16'd5571: out <= 16'hFF76;
    16'd5572: out <= 16'hFFCE;    16'd5573: out <= 16'h036D;    16'd5574: out <= 16'h0088;    16'd5575: out <= 16'hFB3F;
    16'd5576: out <= 16'hFE41;    16'd5577: out <= 16'h057E;    16'd5578: out <= 16'h002D;    16'd5579: out <= 16'h0074;
    16'd5580: out <= 16'h0339;    16'd5581: out <= 16'hFA4E;    16'd5582: out <= 16'hF747;    16'd5583: out <= 16'h03B8;
    16'd5584: out <= 16'hFE5E;    16'd5585: out <= 16'hFC7F;    16'd5586: out <= 16'hFD64;    16'd5587: out <= 16'h04E2;
    16'd5588: out <= 16'h028C;    16'd5589: out <= 16'h010E;    16'd5590: out <= 16'h0678;    16'd5591: out <= 16'h03C4;
    16'd5592: out <= 16'hFDCF;    16'd5593: out <= 16'h03A5;    16'd5594: out <= 16'hFE3C;    16'd5595: out <= 16'hF930;
    16'd5596: out <= 16'hF8C5;    16'd5597: out <= 16'h0034;    16'd5598: out <= 16'hF978;    16'd5599: out <= 16'hFA90;
    16'd5600: out <= 16'h00E5;    16'd5601: out <= 16'hFF6F;    16'd5602: out <= 16'hFDEB;    16'd5603: out <= 16'hFB7B;
    16'd5604: out <= 16'h02F1;    16'd5605: out <= 16'hFFFC;    16'd5606: out <= 16'hFCBF;    16'd5607: out <= 16'h0510;
    16'd5608: out <= 16'hFCC6;    16'd5609: out <= 16'hFE31;    16'd5610: out <= 16'hF623;    16'd5611: out <= 16'hFF7F;
    16'd5612: out <= 16'h085D;    16'd5613: out <= 16'hFDB5;    16'd5614: out <= 16'hF7AA;    16'd5615: out <= 16'h0171;
    16'd5616: out <= 16'h064E;    16'd5617: out <= 16'h03C0;    16'd5618: out <= 16'h013E;    16'd5619: out <= 16'h00E5;
    16'd5620: out <= 16'h02EE;    16'd5621: out <= 16'hFFF7;    16'd5622: out <= 16'h0296;    16'd5623: out <= 16'h00DB;
    16'd5624: out <= 16'hFB06;    16'd5625: out <= 16'hFAB4;    16'd5626: out <= 16'hFAD3;    16'd5627: out <= 16'h0256;
    16'd5628: out <= 16'hFCED;    16'd5629: out <= 16'hFD17;    16'd5630: out <= 16'h0320;    16'd5631: out <= 16'hFBC4;
    16'd5632: out <= 16'hFB51;    16'd5633: out <= 16'h0041;    16'd5634: out <= 16'h011F;    16'd5635: out <= 16'h049D;
    16'd5636: out <= 16'h0087;    16'd5637: out <= 16'hFF36;    16'd5638: out <= 16'h01DD;    16'd5639: out <= 16'hFCA0;
    16'd5640: out <= 16'hF9B1;    16'd5641: out <= 16'h039F;    16'd5642: out <= 16'h02DB;    16'd5643: out <= 16'hFD11;
    16'd5644: out <= 16'hFE4B;    16'd5645: out <= 16'h0383;    16'd5646: out <= 16'hFCCD;    16'd5647: out <= 16'hFC63;
    16'd5648: out <= 16'hF611;    16'd5649: out <= 16'hFE50;    16'd5650: out <= 16'h0274;    16'd5651: out <= 16'h0292;
    16'd5652: out <= 16'hFDE4;    16'd5653: out <= 16'h050D;    16'd5654: out <= 16'h072D;    16'd5655: out <= 16'hFA3F;
    16'd5656: out <= 16'hFA99;    16'd5657: out <= 16'hFCFC;    16'd5658: out <= 16'hFE2A;    16'd5659: out <= 16'hFB82;
    16'd5660: out <= 16'h0082;    16'd5661: out <= 16'h002B;    16'd5662: out <= 16'hFE60;    16'd5663: out <= 16'h0675;
    16'd5664: out <= 16'h0089;    16'd5665: out <= 16'hFFEA;    16'd5666: out <= 16'h05AA;    16'd5667: out <= 16'hFD8F;
    16'd5668: out <= 16'h063A;    16'd5669: out <= 16'h0284;    16'd5670: out <= 16'h0015;    16'd5671: out <= 16'h0011;
    16'd5672: out <= 16'h03C2;    16'd5673: out <= 16'h0061;    16'd5674: out <= 16'hF861;    16'd5675: out <= 16'hFBFE;
    16'd5676: out <= 16'h01E7;    16'd5677: out <= 16'h003D;    16'd5678: out <= 16'hFC87;    16'd5679: out <= 16'h0168;
    16'd5680: out <= 16'hFA8E;    16'd5681: out <= 16'hFD6E;    16'd5682: out <= 16'hFD02;    16'd5683: out <= 16'h0488;
    16'd5684: out <= 16'h02DC;    16'd5685: out <= 16'hFBDE;    16'd5686: out <= 16'h02E1;    16'd5687: out <= 16'h034F;
    16'd5688: out <= 16'h09E2;    16'd5689: out <= 16'h01B4;    16'd5690: out <= 16'h0379;    16'd5691: out <= 16'h03D8;
    16'd5692: out <= 16'hFFFC;    16'd5693: out <= 16'hFF3E;    16'd5694: out <= 16'h0396;    16'd5695: out <= 16'h060B;
    16'd5696: out <= 16'h0D2B;    16'd5697: out <= 16'h03E2;    16'd5698: out <= 16'h03B7;    16'd5699: out <= 16'h043A;
    16'd5700: out <= 16'h0532;    16'd5701: out <= 16'hFD7B;    16'd5702: out <= 16'h022D;    16'd5703: out <= 16'h002E;
    16'd5704: out <= 16'h0667;    16'd5705: out <= 16'hFE9F;    16'd5706: out <= 16'h032A;    16'd5707: out <= 16'h0387;
    16'd5708: out <= 16'h0558;    16'd5709: out <= 16'h03C7;    16'd5710: out <= 16'h078C;    16'd5711: out <= 16'h08D8;
    16'd5712: out <= 16'h0848;    16'd5713: out <= 16'h050F;    16'd5714: out <= 16'h07E7;    16'd5715: out <= 16'h056C;
    16'd5716: out <= 16'h00C3;    16'd5717: out <= 16'h03A8;    16'd5718: out <= 16'h0A1B;    16'd5719: out <= 16'hFF75;
    16'd5720: out <= 16'h035D;    16'd5721: out <= 16'hF8CB;    16'd5722: out <= 16'h07EF;    16'd5723: out <= 16'hFD71;
    16'd5724: out <= 16'h01EE;    16'd5725: out <= 16'h05F0;    16'd5726: out <= 16'h05BB;    16'd5727: out <= 16'h0808;
    16'd5728: out <= 16'h038D;    16'd5729: out <= 16'h02FF;    16'd5730: out <= 16'h046A;    16'd5731: out <= 16'h0119;
    16'd5732: out <= 16'h0717;    16'd5733: out <= 16'h0421;    16'd5734: out <= 16'h0527;    16'd5735: out <= 16'h07AA;
    16'd5736: out <= 16'h09C4;    16'd5737: out <= 16'hFE6B;    16'd5738: out <= 16'h0504;    16'd5739: out <= 16'h01C8;
    16'd5740: out <= 16'h0189;    16'd5741: out <= 16'h030F;    16'd5742: out <= 16'h017B;    16'd5743: out <= 16'hFE44;
    16'd5744: out <= 16'h015B;    16'd5745: out <= 16'h04DF;    16'd5746: out <= 16'h0678;    16'd5747: out <= 16'h058C;
    16'd5748: out <= 16'h050D;    16'd5749: out <= 16'h0297;    16'd5750: out <= 16'hFFAC;    16'd5751: out <= 16'h042F;
    16'd5752: out <= 16'hFDC9;    16'd5753: out <= 16'h0626;    16'd5754: out <= 16'h0347;    16'd5755: out <= 16'h0280;
    16'd5756: out <= 16'h07A0;    16'd5757: out <= 16'h03F3;    16'd5758: out <= 16'h024C;    16'd5759: out <= 16'h06B1;
    16'd5760: out <= 16'hFD48;    16'd5761: out <= 16'h03B4;    16'd5762: out <= 16'h03C1;    16'd5763: out <= 16'h02E5;
    16'd5764: out <= 16'h062B;    16'd5765: out <= 16'h0E28;    16'd5766: out <= 16'h02A5;    16'd5767: out <= 16'h05DE;
    16'd5768: out <= 16'h0B60;    16'd5769: out <= 16'h0751;    16'd5770: out <= 16'h054A;    16'd5771: out <= 16'hF8D3;
    16'd5772: out <= 16'h0A03;    16'd5773: out <= 16'h0567;    16'd5774: out <= 16'h0076;    16'd5775: out <= 16'hFDEC;
    16'd5776: out <= 16'h0698;    16'd5777: out <= 16'h0625;    16'd5778: out <= 16'h0441;    16'd5779: out <= 16'hFD7F;
    16'd5780: out <= 16'h04E9;    16'd5781: out <= 16'h03ED;    16'd5782: out <= 16'h08F2;    16'd5783: out <= 16'hFF87;
    16'd5784: out <= 16'h00DC;    16'd5785: out <= 16'hFF74;    16'd5786: out <= 16'h06D4;    16'd5787: out <= 16'h01C9;
    16'd5788: out <= 16'h05D4;    16'd5789: out <= 16'h06A9;    16'd5790: out <= 16'h0A7D;    16'd5791: out <= 16'h0CA0;
    16'd5792: out <= 16'h0A35;    16'd5793: out <= 16'h027A;    16'd5794: out <= 16'h05AC;    16'd5795: out <= 16'h0354;
    16'd5796: out <= 16'h0BCE;    16'd5797: out <= 16'hFE76;    16'd5798: out <= 16'h0375;    16'd5799: out <= 16'hFDC3;
    16'd5800: out <= 16'h09DD;    16'd5801: out <= 16'h0A6C;    16'd5802: out <= 16'h06EC;    16'd5803: out <= 16'h0222;
    16'd5804: out <= 16'h04A2;    16'd5805: out <= 16'h016C;    16'd5806: out <= 16'h054A;    16'd5807: out <= 16'h05C9;
    16'd5808: out <= 16'h04F4;    16'd5809: out <= 16'h01CD;    16'd5810: out <= 16'h00B5;    16'd5811: out <= 16'h017D;
    16'd5812: out <= 16'h009E;    16'd5813: out <= 16'h0863;    16'd5814: out <= 16'h023B;    16'd5815: out <= 16'h082C;
    16'd5816: out <= 16'h059B;    16'd5817: out <= 16'h03B4;    16'd5818: out <= 16'h06A9;    16'd5819: out <= 16'hFFBD;
    16'd5820: out <= 16'h0759;    16'd5821: out <= 16'h0567;    16'd5822: out <= 16'h0375;    16'd5823: out <= 16'h0333;
    16'd5824: out <= 16'hFD7B;    16'd5825: out <= 16'h02DA;    16'd5826: out <= 16'hFE34;    16'd5827: out <= 16'hFB1B;
    16'd5828: out <= 16'hFE25;    16'd5829: out <= 16'h00BE;    16'd5830: out <= 16'hFE4A;    16'd5831: out <= 16'hFDE0;
    16'd5832: out <= 16'hFEDC;    16'd5833: out <= 16'hFDB6;    16'd5834: out <= 16'h027F;    16'd5835: out <= 16'h0419;
    16'd5836: out <= 16'h04BB;    16'd5837: out <= 16'h02F8;    16'd5838: out <= 16'h004E;    16'd5839: out <= 16'hFE58;
    16'd5840: out <= 16'hFF1C;    16'd5841: out <= 16'h0112;    16'd5842: out <= 16'h0368;    16'd5843: out <= 16'h01DB;
    16'd5844: out <= 16'h0614;    16'd5845: out <= 16'hFFA9;    16'd5846: out <= 16'hFCCB;    16'd5847: out <= 16'hFF68;
    16'd5848: out <= 16'hFEB0;    16'd5849: out <= 16'hFB53;    16'd5850: out <= 16'h0105;    16'd5851: out <= 16'h07DD;
    16'd5852: out <= 16'hF9D1;    16'd5853: out <= 16'hFD74;    16'd5854: out <= 16'h05CF;    16'd5855: out <= 16'h05AD;
    16'd5856: out <= 16'hFF2B;    16'd5857: out <= 16'h0149;    16'd5858: out <= 16'hFEE8;    16'd5859: out <= 16'h01E4;
    16'd5860: out <= 16'hF9D0;    16'd5861: out <= 16'h027F;    16'd5862: out <= 16'hFE8E;    16'd5863: out <= 16'hFE48;
    16'd5864: out <= 16'hFCC7;    16'd5865: out <= 16'hFE0C;    16'd5866: out <= 16'h064D;    16'd5867: out <= 16'hFF1B;
    16'd5868: out <= 16'hF3C1;    16'd5869: out <= 16'hF994;    16'd5870: out <= 16'hFD70;    16'd5871: out <= 16'hFF7B;
    16'd5872: out <= 16'h02B1;    16'd5873: out <= 16'h0308;    16'd5874: out <= 16'hFC76;    16'd5875: out <= 16'hF23A;
    16'd5876: out <= 16'hFCF0;    16'd5877: out <= 16'hF4E9;    16'd5878: out <= 16'h03C2;    16'd5879: out <= 16'hFBEC;
    16'd5880: out <= 16'h013C;    16'd5881: out <= 16'h08A8;    16'd5882: out <= 16'h01FC;    16'd5883: out <= 16'h0167;
    16'd5884: out <= 16'h04C3;    16'd5885: out <= 16'h02E7;    16'd5886: out <= 16'h0000;    16'd5887: out <= 16'h03A1;
    16'd5888: out <= 16'hFAA8;    16'd5889: out <= 16'hFD05;    16'd5890: out <= 16'h073E;    16'd5891: out <= 16'hFC07;
    16'd5892: out <= 16'h091F;    16'd5893: out <= 16'h01E3;    16'd5894: out <= 16'h000F;    16'd5895: out <= 16'hF7EF;
    16'd5896: out <= 16'hF9D5;    16'd5897: out <= 16'hFE8A;    16'd5898: out <= 16'hFD49;    16'd5899: out <= 16'hFC50;
    16'd5900: out <= 16'hF7CB;    16'd5901: out <= 16'hFFD6;    16'd5902: out <= 16'h006A;    16'd5903: out <= 16'hFE2D;
    16'd5904: out <= 16'hFCDF;    16'd5905: out <= 16'h0282;    16'd5906: out <= 16'hFC0A;    16'd5907: out <= 16'hFB18;
    16'd5908: out <= 16'hFA07;    16'd5909: out <= 16'h0327;    16'd5910: out <= 16'hFE40;    16'd5911: out <= 16'h025D;
    16'd5912: out <= 16'hFDE4;    16'd5913: out <= 16'h0235;    16'd5914: out <= 16'hFC1B;    16'd5915: out <= 16'hFDEB;
    16'd5916: out <= 16'h0295;    16'd5917: out <= 16'h0130;    16'd5918: out <= 16'h04AA;    16'd5919: out <= 16'h02E7;
    16'd5920: out <= 16'h0426;    16'd5921: out <= 16'h0C17;    16'd5922: out <= 16'h019B;    16'd5923: out <= 16'hFB09;
    16'd5924: out <= 16'h018B;    16'd5925: out <= 16'h016C;    16'd5926: out <= 16'hFAE7;    16'd5927: out <= 16'h0644;
    16'd5928: out <= 16'hFC00;    16'd5929: out <= 16'hFCB2;    16'd5930: out <= 16'h00DA;    16'd5931: out <= 16'h014B;
    16'd5932: out <= 16'h0358;    16'd5933: out <= 16'h02C1;    16'd5934: out <= 16'hF8F1;    16'd5935: out <= 16'hFDA0;
    16'd5936: out <= 16'hF889;    16'd5937: out <= 16'hFB7B;    16'd5938: out <= 16'hFCB9;    16'd5939: out <= 16'hFDEE;
    16'd5940: out <= 16'h091A;    16'd5941: out <= 16'h02FC;    16'd5942: out <= 16'hFF2D;    16'd5943: out <= 16'h0854;
    16'd5944: out <= 16'h0336;    16'd5945: out <= 16'h0CB5;    16'd5946: out <= 16'h01F0;    16'd5947: out <= 16'h0049;
    16'd5948: out <= 16'hFE41;    16'd5949: out <= 16'h0BAA;    16'd5950: out <= 16'h0BBF;    16'd5951: out <= 16'hFF7E;
    16'd5952: out <= 16'hFFE5;    16'd5953: out <= 16'h0741;    16'd5954: out <= 16'h05F1;    16'd5955: out <= 16'hFECE;
    16'd5956: out <= 16'hFF76;    16'd5957: out <= 16'h001A;    16'd5958: out <= 16'h0261;    16'd5959: out <= 16'h0378;
    16'd5960: out <= 16'h000C;    16'd5961: out <= 16'h038B;    16'd5962: out <= 16'h00B3;    16'd5963: out <= 16'h015F;
    16'd5964: out <= 16'h0446;    16'd5965: out <= 16'h0A9E;    16'd5966: out <= 16'h02B0;    16'd5967: out <= 16'h047D;
    16'd5968: out <= 16'h00D1;    16'd5969: out <= 16'h0530;    16'd5970: out <= 16'h0355;    16'd5971: out <= 16'h039D;
    16'd5972: out <= 16'h017E;    16'd5973: out <= 16'h01D0;    16'd5974: out <= 16'h05EA;    16'd5975: out <= 16'hFEA0;
    16'd5976: out <= 16'h0178;    16'd5977: out <= 16'hFC4D;    16'd5978: out <= 16'h0124;    16'd5979: out <= 16'h06D7;
    16'd5980: out <= 16'h0145;    16'd5981: out <= 16'h032F;    16'd5982: out <= 16'h0985;    16'd5983: out <= 16'h0604;
    16'd5984: out <= 16'h0348;    16'd5985: out <= 16'h00FA;    16'd5986: out <= 16'h05A6;    16'd5987: out <= 16'h0E22;
    16'd5988: out <= 16'h0191;    16'd5989: out <= 16'hFCBA;    16'd5990: out <= 16'h0811;    16'd5991: out <= 16'h0397;
    16'd5992: out <= 16'h02F0;    16'd5993: out <= 16'h0626;    16'd5994: out <= 16'h0137;    16'd5995: out <= 16'h0501;
    16'd5996: out <= 16'h0527;    16'd5997: out <= 16'h021D;    16'd5998: out <= 16'h0026;    16'd5999: out <= 16'h0258;
    16'd6000: out <= 16'h08FF;    16'd6001: out <= 16'h0718;    16'd6002: out <= 16'h0691;    16'd6003: out <= 16'h0709;
    16'd6004: out <= 16'h0451;    16'd6005: out <= 16'h00BE;    16'd6006: out <= 16'hFEB0;    16'd6007: out <= 16'h03FF;
    16'd6008: out <= 16'h09C5;    16'd6009: out <= 16'h0D1A;    16'd6010: out <= 16'hFDAD;    16'd6011: out <= 16'h02F3;
    16'd6012: out <= 16'hFF44;    16'd6013: out <= 16'hFDE6;    16'd6014: out <= 16'h0CBA;    16'd6015: out <= 16'h06E6;
    16'd6016: out <= 16'hFF85;    16'd6017: out <= 16'hFD46;    16'd6018: out <= 16'h0504;    16'd6019: out <= 16'h01E6;
    16'd6020: out <= 16'h05E5;    16'd6021: out <= 16'h0246;    16'd6022: out <= 16'hFE94;    16'd6023: out <= 16'h0741;
    16'd6024: out <= 16'h0962;    16'd6025: out <= 16'h03AC;    16'd6026: out <= 16'h011A;    16'd6027: out <= 16'h06F9;
    16'd6028: out <= 16'h027D;    16'd6029: out <= 16'h048B;    16'd6030: out <= 16'h0678;    16'd6031: out <= 16'h0505;
    16'd6032: out <= 16'h04B5;    16'd6033: out <= 16'hFF5D;    16'd6034: out <= 16'h02CB;    16'd6035: out <= 16'h0349;
    16'd6036: out <= 16'h03CF;    16'd6037: out <= 16'h054D;    16'd6038: out <= 16'hFC84;    16'd6039: out <= 16'h02DF;
    16'd6040: out <= 16'h074D;    16'd6041: out <= 16'h0966;    16'd6042: out <= 16'h0BEA;    16'd6043: out <= 16'h05C5;
    16'd6044: out <= 16'h0813;    16'd6045: out <= 16'h0D59;    16'd6046: out <= 16'h0504;    16'd6047: out <= 16'h069C;
    16'd6048: out <= 16'h01AE;    16'd6049: out <= 16'hFED8;    16'd6050: out <= 16'h0277;    16'd6051: out <= 16'h01F9;
    16'd6052: out <= 16'h070D;    16'd6053: out <= 16'h0127;    16'd6054: out <= 16'h0814;    16'd6055: out <= 16'hFDBB;
    16'd6056: out <= 16'h0371;    16'd6057: out <= 16'h0721;    16'd6058: out <= 16'h00E8;    16'd6059: out <= 16'h06C7;
    16'd6060: out <= 16'h0596;    16'd6061: out <= 16'h06E5;    16'd6062: out <= 16'hFF95;    16'd6063: out <= 16'h03ED;
    16'd6064: out <= 16'hFEA0;    16'd6065: out <= 16'h042C;    16'd6066: out <= 16'h0755;    16'd6067: out <= 16'h060A;
    16'd6068: out <= 16'hFED2;    16'd6069: out <= 16'h0979;    16'd6070: out <= 16'h09AB;    16'd6071: out <= 16'h0418;
    16'd6072: out <= 16'h01C3;    16'd6073: out <= 16'h0161;    16'd6074: out <= 16'h0390;    16'd6075: out <= 16'h063E;
    16'd6076: out <= 16'h05EA;    16'd6077: out <= 16'h0510;    16'd6078: out <= 16'h0127;    16'd6079: out <= 16'h0248;
    16'd6080: out <= 16'h0502;    16'd6081: out <= 16'hFE51;    16'd6082: out <= 16'hFA54;    16'd6083: out <= 16'h0013;
    16'd6084: out <= 16'h02C0;    16'd6085: out <= 16'h01A0;    16'd6086: out <= 16'hFCBB;    16'd6087: out <= 16'hFE08;
    16'd6088: out <= 16'hFE4D;    16'd6089: out <= 16'h04FA;    16'd6090: out <= 16'h04AB;    16'd6091: out <= 16'hF866;
    16'd6092: out <= 16'h01CA;    16'd6093: out <= 16'hFF8D;    16'd6094: out <= 16'h0176;    16'd6095: out <= 16'h03A4;
    16'd6096: out <= 16'hF7CB;    16'd6097: out <= 16'hFBCD;    16'd6098: out <= 16'h047D;    16'd6099: out <= 16'hFC77;
    16'd6100: out <= 16'h03E9;    16'd6101: out <= 16'h029F;    16'd6102: out <= 16'h0129;    16'd6103: out <= 16'h06F3;
    16'd6104: out <= 16'hF915;    16'd6105: out <= 16'h0CDA;    16'd6106: out <= 16'h02F0;    16'd6107: out <= 16'h0183;
    16'd6108: out <= 16'hFBC4;    16'd6109: out <= 16'h0119;    16'd6110: out <= 16'h007C;    16'd6111: out <= 16'hFBDB;
    16'd6112: out <= 16'hFC1E;    16'd6113: out <= 16'h04AE;    16'd6114: out <= 16'h0007;    16'd6115: out <= 16'hFDDA;
    16'd6116: out <= 16'hF6E7;    16'd6117: out <= 16'h00D6;    16'd6118: out <= 16'h02D1;    16'd6119: out <= 16'h0551;
    16'd6120: out <= 16'hFEB8;    16'd6121: out <= 16'hFABF;    16'd6122: out <= 16'h00C3;    16'd6123: out <= 16'hF8DB;
    16'd6124: out <= 16'hF618;    16'd6125: out <= 16'hFB8A;    16'd6126: out <= 16'hFDEF;    16'd6127: out <= 16'hFDC7;
    16'd6128: out <= 16'h03FE;    16'd6129: out <= 16'hFC88;    16'd6130: out <= 16'h00CA;    16'd6131: out <= 16'h0379;
    16'd6132: out <= 16'hFCFB;    16'd6133: out <= 16'h00BF;    16'd6134: out <= 16'h01F2;    16'd6135: out <= 16'hFCAF;
    16'd6136: out <= 16'hFF2A;    16'd6137: out <= 16'hF73A;    16'd6138: out <= 16'h0366;    16'd6139: out <= 16'hFF2F;
    16'd6140: out <= 16'h01C8;    16'd6141: out <= 16'hF7BF;    16'd6142: out <= 16'h0324;    16'd6143: out <= 16'h03D1;
    16'd6144: out <= 16'hFB2D;    16'd6145: out <= 16'hFF1E;    16'd6146: out <= 16'h05DA;    16'd6147: out <= 16'hFEF5;
    16'd6148: out <= 16'hFE98;    16'd6149: out <= 16'h02A0;    16'd6150: out <= 16'hF7F7;    16'd6151: out <= 16'h0941;
    16'd6152: out <= 16'h00BF;    16'd6153: out <= 16'hFE6D;    16'd6154: out <= 16'hFDD2;    16'd6155: out <= 16'h0519;
    16'd6156: out <= 16'h03FE;    16'd6157: out <= 16'h0155;    16'd6158: out <= 16'h0004;    16'd6159: out <= 16'h0151;
    16'd6160: out <= 16'h0096;    16'd6161: out <= 16'h00E7;    16'd6162: out <= 16'h021E;    16'd6163: out <= 16'hFCA2;
    16'd6164: out <= 16'hFB2A;    16'd6165: out <= 16'hFE75;    16'd6166: out <= 16'hF491;    16'd6167: out <= 16'h012B;
    16'd6168: out <= 16'h014C;    16'd6169: out <= 16'hFD02;    16'd6170: out <= 16'h0375;    16'd6171: out <= 16'hFF3A;
    16'd6172: out <= 16'h052F;    16'd6173: out <= 16'h000D;    16'd6174: out <= 16'hFF9E;    16'd6175: out <= 16'hFF76;
    16'd6176: out <= 16'h0784;    16'd6177: out <= 16'h00E3;    16'd6178: out <= 16'hFC28;    16'd6179: out <= 16'h06BB;
    16'd6180: out <= 16'h07B6;    16'd6181: out <= 16'hF5A0;    16'd6182: out <= 16'hFF4C;    16'd6183: out <= 16'h0411;
    16'd6184: out <= 16'hFF4B;    16'd6185: out <= 16'h0093;    16'd6186: out <= 16'h000C;    16'd6187: out <= 16'h0214;
    16'd6188: out <= 16'h05E4;    16'd6189: out <= 16'hFF1E;    16'd6190: out <= 16'h0487;    16'd6191: out <= 16'hFD03;
    16'd6192: out <= 16'hFAB9;    16'd6193: out <= 16'h0761;    16'd6194: out <= 16'h02CA;    16'd6195: out <= 16'h046A;
    16'd6196: out <= 16'hFEAB;    16'd6197: out <= 16'h058C;    16'd6198: out <= 16'h0B77;    16'd6199: out <= 16'h0692;
    16'd6200: out <= 16'h02C1;    16'd6201: out <= 16'h05A0;    16'd6202: out <= 16'h0161;    16'd6203: out <= 16'h0D84;
    16'd6204: out <= 16'hFF72;    16'd6205: out <= 16'hFA63;    16'd6206: out <= 16'h0225;    16'd6207: out <= 16'h0215;
    16'd6208: out <= 16'h01D8;    16'd6209: out <= 16'h00D4;    16'd6210: out <= 16'h0202;    16'd6211: out <= 16'h02E6;
    16'd6212: out <= 16'h0571;    16'd6213: out <= 16'h0499;    16'd6214: out <= 16'h050E;    16'd6215: out <= 16'h058A;
    16'd6216: out <= 16'h06CA;    16'd6217: out <= 16'hFCE6;    16'd6218: out <= 16'h053E;    16'd6219: out <= 16'h09BD;
    16'd6220: out <= 16'h00CB;    16'd6221: out <= 16'h0284;    16'd6222: out <= 16'h0685;    16'd6223: out <= 16'h0A08;
    16'd6224: out <= 16'h02C9;    16'd6225: out <= 16'h062C;    16'd6226: out <= 16'h09A5;    16'd6227: out <= 16'h0787;
    16'd6228: out <= 16'h029C;    16'd6229: out <= 16'h060C;    16'd6230: out <= 16'h0515;    16'd6231: out <= 16'h024D;
    16'd6232: out <= 16'hFD86;    16'd6233: out <= 16'h0894;    16'd6234: out <= 16'h02BE;    16'd6235: out <= 16'hFE83;
    16'd6236: out <= 16'h0717;    16'd6237: out <= 16'hFE93;    16'd6238: out <= 16'h06E1;    16'd6239: out <= 16'hFEC9;
    16'd6240: out <= 16'h001F;    16'd6241: out <= 16'h02EB;    16'd6242: out <= 16'h0AF1;    16'd6243: out <= 16'h043B;
    16'd6244: out <= 16'h09C0;    16'd6245: out <= 16'h0A4E;    16'd6246: out <= 16'h044D;    16'd6247: out <= 16'h0451;
    16'd6248: out <= 16'h0459;    16'd6249: out <= 16'h0081;    16'd6250: out <= 16'h052F;    16'd6251: out <= 16'h0BC2;
    16'd6252: out <= 16'h0504;    16'd6253: out <= 16'h0255;    16'd6254: out <= 16'h045C;    16'd6255: out <= 16'h02A2;
    16'd6256: out <= 16'h0972;    16'd6257: out <= 16'hFFE7;    16'd6258: out <= 16'h037D;    16'd6259: out <= 16'h04A3;
    16'd6260: out <= 16'hFEA4;    16'd6261: out <= 16'h04AE;    16'd6262: out <= 16'h0496;    16'd6263: out <= 16'h0561;
    16'd6264: out <= 16'hFF5E;    16'd6265: out <= 16'h073A;    16'd6266: out <= 16'h0654;    16'd6267: out <= 16'h05C6;
    16'd6268: out <= 16'h0296;    16'd6269: out <= 16'h02B2;    16'd6270: out <= 16'h0452;    16'd6271: out <= 16'h0A8C;
    16'd6272: out <= 16'h01BA;    16'd6273: out <= 16'h0A0C;    16'd6274: out <= 16'h05A1;    16'd6275: out <= 16'h0347;
    16'd6276: out <= 16'h055D;    16'd6277: out <= 16'h06A0;    16'd6278: out <= 16'h021B;    16'd6279: out <= 16'h0431;
    16'd6280: out <= 16'hFD29;    16'd6281: out <= 16'h03C5;    16'd6282: out <= 16'h0502;    16'd6283: out <= 16'h05E9;
    16'd6284: out <= 16'h0249;    16'd6285: out <= 16'hFECC;    16'd6286: out <= 16'h039E;    16'd6287: out <= 16'h07D9;
    16'd6288: out <= 16'h01B3;    16'd6289: out <= 16'h048B;    16'd6290: out <= 16'h0333;    16'd6291: out <= 16'h0BC8;
    16'd6292: out <= 16'h0369;    16'd6293: out <= 16'h064D;    16'd6294: out <= 16'h0951;    16'd6295: out <= 16'hFF2B;
    16'd6296: out <= 16'h0597;    16'd6297: out <= 16'h00C2;    16'd6298: out <= 16'h052B;    16'd6299: out <= 16'h0013;
    16'd6300: out <= 16'h0C65;    16'd6301: out <= 16'h0250;    16'd6302: out <= 16'h052D;    16'd6303: out <= 16'h0960;
    16'd6304: out <= 16'h070C;    16'd6305: out <= 16'h025D;    16'd6306: out <= 16'h0647;    16'd6307: out <= 16'hFEED;
    16'd6308: out <= 16'h00AE;    16'd6309: out <= 16'h0025;    16'd6310: out <= 16'h0A32;    16'd6311: out <= 16'h012C;
    16'd6312: out <= 16'h0116;    16'd6313: out <= 16'h07C6;    16'd6314: out <= 16'h09AC;    16'd6315: out <= 16'h0E5E;
    16'd6316: out <= 16'h0182;    16'd6317: out <= 16'hFE24;    16'd6318: out <= 16'h0561;    16'd6319: out <= 16'h027B;
    16'd6320: out <= 16'h0466;    16'd6321: out <= 16'h020F;    16'd6322: out <= 16'h0663;    16'd6323: out <= 16'h016A;
    16'd6324: out <= 16'hFE37;    16'd6325: out <= 16'h0BD7;    16'd6326: out <= 16'h02F0;    16'd6327: out <= 16'h007E;
    16'd6328: out <= 16'h0865;    16'd6329: out <= 16'h0209;    16'd6330: out <= 16'h07AE;    16'd6331: out <= 16'h039E;
    16'd6332: out <= 16'h00A0;    16'd6333: out <= 16'h00DF;    16'd6334: out <= 16'h047E;    16'd6335: out <= 16'h09C5;
    16'd6336: out <= 16'h0824;    16'd6337: out <= 16'h064E;    16'd6338: out <= 16'hFA99;    16'd6339: out <= 16'hFFB1;
    16'd6340: out <= 16'hFB87;    16'd6341: out <= 16'hFB87;    16'd6342: out <= 16'h05B8;    16'd6343: out <= 16'h003C;
    16'd6344: out <= 16'h01A2;    16'd6345: out <= 16'h00FF;    16'd6346: out <= 16'hFC78;    16'd6347: out <= 16'hFCBE;
    16'd6348: out <= 16'h03C7;    16'd6349: out <= 16'h00D8;    16'd6350: out <= 16'hFECC;    16'd6351: out <= 16'h0111;
    16'd6352: out <= 16'hFB40;    16'd6353: out <= 16'hFE23;    16'd6354: out <= 16'hF864;    16'd6355: out <= 16'h09F6;
    16'd6356: out <= 16'h034C;    16'd6357: out <= 16'h05E3;    16'd6358: out <= 16'h010D;    16'd6359: out <= 16'h00BD;
    16'd6360: out <= 16'h00DB;    16'd6361: out <= 16'hFC93;    16'd6362: out <= 16'hF5FF;    16'd6363: out <= 16'h0028;
    16'd6364: out <= 16'hFF83;    16'd6365: out <= 16'hFF5B;    16'd6366: out <= 16'h00B6;    16'd6367: out <= 16'hFC59;
    16'd6368: out <= 16'hFC1D;    16'd6369: out <= 16'hFFD1;    16'd6370: out <= 16'hF6EE;    16'd6371: out <= 16'hFC84;
    16'd6372: out <= 16'h015A;    16'd6373: out <= 16'hFA80;    16'd6374: out <= 16'h0121;    16'd6375: out <= 16'h016F;
    16'd6376: out <= 16'h01B1;    16'd6377: out <= 16'hFF85;    16'd6378: out <= 16'hFEAF;    16'd6379: out <= 16'h0981;
    16'd6380: out <= 16'h012D;    16'd6381: out <= 16'hFC81;    16'd6382: out <= 16'hFCC7;    16'd6383: out <= 16'hFF62;
    16'd6384: out <= 16'h01AA;    16'd6385: out <= 16'hFDC4;    16'd6386: out <= 16'h0064;    16'd6387: out <= 16'h028E;
    16'd6388: out <= 16'hFBE7;    16'd6389: out <= 16'hFF43;    16'd6390: out <= 16'h05DD;    16'd6391: out <= 16'h0225;
    16'd6392: out <= 16'h03A7;    16'd6393: out <= 16'hFE15;    16'd6394: out <= 16'h032F;    16'd6395: out <= 16'hFC4F;
    16'd6396: out <= 16'hFEC1;    16'd6397: out <= 16'h0387;    16'd6398: out <= 16'h02DB;    16'd6399: out <= 16'h0240;
    16'd6400: out <= 16'hFD74;    16'd6401: out <= 16'hFEE8;    16'd6402: out <= 16'hFE01;    16'd6403: out <= 16'h0197;
    16'd6404: out <= 16'hF9AD;    16'd6405: out <= 16'h0712;    16'd6406: out <= 16'hFB56;    16'd6407: out <= 16'h02DF;
    16'd6408: out <= 16'hFDC8;    16'd6409: out <= 16'hFE43;    16'd6410: out <= 16'hFEBE;    16'd6411: out <= 16'hFEF0;
    16'd6412: out <= 16'hFCC1;    16'd6413: out <= 16'hFC77;    16'd6414: out <= 16'hFEC6;    16'd6415: out <= 16'h0062;
    16'd6416: out <= 16'hFC79;    16'd6417: out <= 16'hFE95;    16'd6418: out <= 16'h00B3;    16'd6419: out <= 16'hF833;
    16'd6420: out <= 16'h006D;    16'd6421: out <= 16'h00E4;    16'd6422: out <= 16'h0086;    16'd6423: out <= 16'hF918;
    16'd6424: out <= 16'h00B2;    16'd6425: out <= 16'hFFDE;    16'd6426: out <= 16'h024B;    16'd6427: out <= 16'h0009;
    16'd6428: out <= 16'hFAE0;    16'd6429: out <= 16'hF827;    16'd6430: out <= 16'h0643;    16'd6431: out <= 16'h01AA;
    16'd6432: out <= 16'hFB1E;    16'd6433: out <= 16'hF8D6;    16'd6434: out <= 16'h00D5;    16'd6435: out <= 16'h03AD;
    16'd6436: out <= 16'hFE6C;    16'd6437: out <= 16'hFCD1;    16'd6438: out <= 16'hFE77;    16'd6439: out <= 16'h004E;
    16'd6440: out <= 16'h0038;    16'd6441: out <= 16'hFDA6;    16'd6442: out <= 16'h0098;    16'd6443: out <= 16'hF8F3;
    16'd6444: out <= 16'h0140;    16'd6445: out <= 16'hFD70;    16'd6446: out <= 16'hFD78;    16'd6447: out <= 16'hFFA5;
    16'd6448: out <= 16'hFE4C;    16'd6449: out <= 16'hFCB5;    16'd6450: out <= 16'h084F;    16'd6451: out <= 16'h04BB;
    16'd6452: out <= 16'h0464;    16'd6453: out <= 16'h00D0;    16'd6454: out <= 16'h03B4;    16'd6455: out <= 16'h086C;
    16'd6456: out <= 16'h065A;    16'd6457: out <= 16'h039F;    16'd6458: out <= 16'hFE2E;    16'd6459: out <= 16'h07DB;
    16'd6460: out <= 16'h04CD;    16'd6461: out <= 16'h0413;    16'd6462: out <= 16'h0324;    16'd6463: out <= 16'hFD72;
    16'd6464: out <= 16'h0332;    16'd6465: out <= 16'h0781;    16'd6466: out <= 16'h07B1;    16'd6467: out <= 16'h0334;
    16'd6468: out <= 16'h09C4;    16'd6469: out <= 16'h0376;    16'd6470: out <= 16'h09D4;    16'd6471: out <= 16'h060E;
    16'd6472: out <= 16'h044E;    16'd6473: out <= 16'h0D3C;    16'd6474: out <= 16'h0330;    16'd6475: out <= 16'h0C9D;
    16'd6476: out <= 16'h0942;    16'd6477: out <= 16'hFF06;    16'd6478: out <= 16'h080A;    16'd6479: out <= 16'h0614;
    16'd6480: out <= 16'hFF2C;    16'd6481: out <= 16'h03DF;    16'd6482: out <= 16'h09DE;    16'd6483: out <= 16'h07B3;
    16'd6484: out <= 16'h0A6A;    16'd6485: out <= 16'h0C01;    16'd6486: out <= 16'h0ACD;    16'd6487: out <= 16'hFC83;
    16'd6488: out <= 16'h048C;    16'd6489: out <= 16'h04F8;    16'd6490: out <= 16'h0795;    16'd6491: out <= 16'h0B9C;
    16'd6492: out <= 16'h0498;    16'd6493: out <= 16'h0682;    16'd6494: out <= 16'h052E;    16'd6495: out <= 16'h0204;
    16'd6496: out <= 16'hFF35;    16'd6497: out <= 16'hFD5F;    16'd6498: out <= 16'h0150;    16'd6499: out <= 16'h0661;
    16'd6500: out <= 16'h03EB;    16'd6501: out <= 16'h0308;    16'd6502: out <= 16'h0321;    16'd6503: out <= 16'h05EB;
    16'd6504: out <= 16'h0604;    16'd6505: out <= 16'hFE8F;    16'd6506: out <= 16'h0417;    16'd6507: out <= 16'h104E;
    16'd6508: out <= 16'hFF48;    16'd6509: out <= 16'hFBA4;    16'd6510: out <= 16'h08E1;    16'd6511: out <= 16'hFF6F;
    16'd6512: out <= 16'hFFBE;    16'd6513: out <= 16'h072E;    16'd6514: out <= 16'h0662;    16'd6515: out <= 16'h0435;
    16'd6516: out <= 16'h0995;    16'd6517: out <= 16'h0A42;    16'd6518: out <= 16'h0C0A;    16'd6519: out <= 16'h0487;
    16'd6520: out <= 16'h06B7;    16'd6521: out <= 16'h04F9;    16'd6522: out <= 16'h00D9;    16'd6523: out <= 16'h0196;
    16'd6524: out <= 16'h0506;    16'd6525: out <= 16'hFAA1;    16'd6526: out <= 16'h072D;    16'd6527: out <= 16'h0526;
    16'd6528: out <= 16'h0813;    16'd6529: out <= 16'h05B2;    16'd6530: out <= 16'h08EA;    16'd6531: out <= 16'h0422;
    16'd6532: out <= 16'hFC74;    16'd6533: out <= 16'h0514;    16'd6534: out <= 16'h016C;    16'd6535: out <= 16'h0641;
    16'd6536: out <= 16'h0275;    16'd6537: out <= 16'hFDBC;    16'd6538: out <= 16'h01D4;    16'd6539: out <= 16'h0574;
    16'd6540: out <= 16'h0104;    16'd6541: out <= 16'h0683;    16'd6542: out <= 16'h0386;    16'd6543: out <= 16'h06D1;
    16'd6544: out <= 16'h0514;    16'd6545: out <= 16'h01F1;    16'd6546: out <= 16'h03DA;    16'd6547: out <= 16'h018B;
    16'd6548: out <= 16'h0912;    16'd6549: out <= 16'h0569;    16'd6550: out <= 16'h03FD;    16'd6551: out <= 16'h03D2;
    16'd6552: out <= 16'h05D3;    16'd6553: out <= 16'h09BB;    16'd6554: out <= 16'h014B;    16'd6555: out <= 16'h0795;
    16'd6556: out <= 16'h02DA;    16'd6557: out <= 16'h0586;    16'd6558: out <= 16'h04A6;    16'd6559: out <= 16'h07F4;
    16'd6560: out <= 16'h0670;    16'd6561: out <= 16'h04DC;    16'd6562: out <= 16'h0178;    16'd6563: out <= 16'h03FB;
    16'd6564: out <= 16'hFD52;    16'd6565: out <= 16'h0C46;    16'd6566: out <= 16'h0A98;    16'd6567: out <= 16'hFE3E;
    16'd6568: out <= 16'h0630;    16'd6569: out <= 16'h031E;    16'd6570: out <= 16'h029C;    16'd6571: out <= 16'h011A;
    16'd6572: out <= 16'h0380;    16'd6573: out <= 16'hFE9D;    16'd6574: out <= 16'h0EF7;    16'd6575: out <= 16'hFC78;
    16'd6576: out <= 16'h0069;    16'd6577: out <= 16'h0A53;    16'd6578: out <= 16'h0304;    16'd6579: out <= 16'h08D3;
    16'd6580: out <= 16'h0375;    16'd6581: out <= 16'h06B0;    16'd6582: out <= 16'h07E4;    16'd6583: out <= 16'h06E8;
    16'd6584: out <= 16'h00E2;    16'd6585: out <= 16'h0C76;    16'd6586: out <= 16'h0670;    16'd6587: out <= 16'h069A;
    16'd6588: out <= 16'h04C4;    16'd6589: out <= 16'h049E;    16'd6590: out <= 16'hFE4B;    16'd6591: out <= 16'hFFB2;
    16'd6592: out <= 16'h00C1;    16'd6593: out <= 16'hFE5C;    16'd6594: out <= 16'h074C;    16'd6595: out <= 16'h0671;
    16'd6596: out <= 16'h0789;    16'd6597: out <= 16'h00C3;    16'd6598: out <= 16'h0195;    16'd6599: out <= 16'hF955;
    16'd6600: out <= 16'hFE61;    16'd6601: out <= 16'h0057;    16'd6602: out <= 16'h003B;    16'd6603: out <= 16'h0292;
    16'd6604: out <= 16'hFBE7;    16'd6605: out <= 16'hFB5F;    16'd6606: out <= 16'hFC1F;    16'd6607: out <= 16'h0403;
    16'd6608: out <= 16'h01EC;    16'd6609: out <= 16'h0687;    16'd6610: out <= 16'hFF50;    16'd6611: out <= 16'hFFEF;
    16'd6612: out <= 16'h051A;    16'd6613: out <= 16'h0256;    16'd6614: out <= 16'h00F9;    16'd6615: out <= 16'hFF91;
    16'd6616: out <= 16'h04AA;    16'd6617: out <= 16'hF9BC;    16'd6618: out <= 16'h030E;    16'd6619: out <= 16'h0712;
    16'd6620: out <= 16'h01B0;    16'd6621: out <= 16'h0697;    16'd6622: out <= 16'h079E;    16'd6623: out <= 16'h023F;
    16'd6624: out <= 16'hFEA7;    16'd6625: out <= 16'h0060;    16'd6626: out <= 16'h026F;    16'd6627: out <= 16'hFE75;
    16'd6628: out <= 16'hFC8E;    16'd6629: out <= 16'hFFBE;    16'd6630: out <= 16'h0339;    16'd6631: out <= 16'hFE80;
    16'd6632: out <= 16'hFE38;    16'd6633: out <= 16'hFCFC;    16'd6634: out <= 16'hF88E;    16'd6635: out <= 16'hFE6C;
    16'd6636: out <= 16'h05F5;    16'd6637: out <= 16'hF82B;    16'd6638: out <= 16'hFCF5;    16'd6639: out <= 16'hFF94;
    16'd6640: out <= 16'hFC8D;    16'd6641: out <= 16'h037F;    16'd6642: out <= 16'h0409;    16'd6643: out <= 16'h04EE;
    16'd6644: out <= 16'h052E;    16'd6645: out <= 16'h0037;    16'd6646: out <= 16'h0B6D;    16'd6647: out <= 16'hFE98;
    16'd6648: out <= 16'hF90E;    16'd6649: out <= 16'hFD06;    16'd6650: out <= 16'h030E;    16'd6651: out <= 16'hFDB3;
    16'd6652: out <= 16'h0136;    16'd6653: out <= 16'hFF77;    16'd6654: out <= 16'hFEA3;    16'd6655: out <= 16'hFF80;
    16'd6656: out <= 16'hF89B;    16'd6657: out <= 16'h00D5;    16'd6658: out <= 16'hFE44;    16'd6659: out <= 16'h0122;
    16'd6660: out <= 16'h003C;    16'd6661: out <= 16'h0025;    16'd6662: out <= 16'hF94A;    16'd6663: out <= 16'hFACA;
    16'd6664: out <= 16'h0132;    16'd6665: out <= 16'h01DC;    16'd6666: out <= 16'hFF20;    16'd6667: out <= 16'hFF01;
    16'd6668: out <= 16'hFE1A;    16'd6669: out <= 16'h00C0;    16'd6670: out <= 16'h006F;    16'd6671: out <= 16'hFCD9;
    16'd6672: out <= 16'h0191;    16'd6673: out <= 16'h0109;    16'd6674: out <= 16'h05F2;    16'd6675: out <= 16'hFF80;
    16'd6676: out <= 16'hFB9D;    16'd6677: out <= 16'hFE64;    16'd6678: out <= 16'hFB95;    16'd6679: out <= 16'h01F1;
    16'd6680: out <= 16'hFAC1;    16'd6681: out <= 16'hFC99;    16'd6682: out <= 16'hFD9C;    16'd6683: out <= 16'h0434;
    16'd6684: out <= 16'h0325;    16'd6685: out <= 16'h01DB;    16'd6686: out <= 16'h01B7;    16'd6687: out <= 16'hFEEF;
    16'd6688: out <= 16'hFED6;    16'd6689: out <= 16'hFB12;    16'd6690: out <= 16'hFD9B;    16'd6691: out <= 16'hFCA2;
    16'd6692: out <= 16'hFA7B;    16'd6693: out <= 16'hFF4B;    16'd6694: out <= 16'hFEE7;    16'd6695: out <= 16'h009F;
    16'd6696: out <= 16'h080A;    16'd6697: out <= 16'hFFCE;    16'd6698: out <= 16'h024B;    16'd6699: out <= 16'hFC1D;
    16'd6700: out <= 16'hF935;    16'd6701: out <= 16'hFB66;    16'd6702: out <= 16'h0136;    16'd6703: out <= 16'h0657;
    16'd6704: out <= 16'hFAE5;    16'd6705: out <= 16'h02E2;    16'd6706: out <= 16'hFFCC;    16'd6707: out <= 16'h0694;
    16'd6708: out <= 16'h002E;    16'd6709: out <= 16'hFFE6;    16'd6710: out <= 16'h00EB;    16'd6711: out <= 16'h0781;
    16'd6712: out <= 16'hFE10;    16'd6713: out <= 16'h0623;    16'd6714: out <= 16'hFECD;    16'd6715: out <= 16'h0887;
    16'd6716: out <= 16'h03F0;    16'd6717: out <= 16'hFADB;    16'd6718: out <= 16'h0604;    16'd6719: out <= 16'h02CF;
    16'd6720: out <= 16'hFB48;    16'd6721: out <= 16'hFECB;    16'd6722: out <= 16'hFE46;    16'd6723: out <= 16'hFEBB;
    16'd6724: out <= 16'h01CF;    16'd6725: out <= 16'h06BE;    16'd6726: out <= 16'h031C;    16'd6727: out <= 16'h0334;
    16'd6728: out <= 16'h0D31;    16'd6729: out <= 16'h03BC;    16'd6730: out <= 16'h0164;    16'd6731: out <= 16'h0CF9;
    16'd6732: out <= 16'h065C;    16'd6733: out <= 16'hFE65;    16'd6734: out <= 16'h08D4;    16'd6735: out <= 16'h05F1;
    16'd6736: out <= 16'h04E1;    16'd6737: out <= 16'h038C;    16'd6738: out <= 16'h000F;    16'd6739: out <= 16'h0290;
    16'd6740: out <= 16'h0678;    16'd6741: out <= 16'h0C35;    16'd6742: out <= 16'h0493;    16'd6743: out <= 16'hFEBA;
    16'd6744: out <= 16'h093A;    16'd6745: out <= 16'h07B5;    16'd6746: out <= 16'h0037;    16'd6747: out <= 16'h074D;
    16'd6748: out <= 16'h07F8;    16'd6749: out <= 16'h087E;    16'd6750: out <= 16'h00E9;    16'd6751: out <= 16'h03B8;
    16'd6752: out <= 16'h0781;    16'd6753: out <= 16'h0255;    16'd6754: out <= 16'h06D0;    16'd6755: out <= 16'h047A;
    16'd6756: out <= 16'h055E;    16'd6757: out <= 16'h0928;    16'd6758: out <= 16'h07A9;    16'd6759: out <= 16'h0510;
    16'd6760: out <= 16'h059F;    16'd6761: out <= 16'h017A;    16'd6762: out <= 16'h0312;    16'd6763: out <= 16'h0279;
    16'd6764: out <= 16'h0781;    16'd6765: out <= 16'h0807;    16'd6766: out <= 16'h0459;    16'd6767: out <= 16'h0104;
    16'd6768: out <= 16'h0265;    16'd6769: out <= 16'h09F1;    16'd6770: out <= 16'h007C;    16'd6771: out <= 16'h0211;
    16'd6772: out <= 16'h07DB;    16'd6773: out <= 16'h0B34;    16'd6774: out <= 16'h0A0C;    16'd6775: out <= 16'h0413;
    16'd6776: out <= 16'h0995;    16'd6777: out <= 16'h0321;    16'd6778: out <= 16'h06A1;    16'd6779: out <= 16'h0699;
    16'd6780: out <= 16'hFF58;    16'd6781: out <= 16'h0549;    16'd6782: out <= 16'h037E;    16'd6783: out <= 16'h0CEC;
    16'd6784: out <= 16'h070E;    16'd6785: out <= 16'h097C;    16'd6786: out <= 16'h00E3;    16'd6787: out <= 16'h0264;
    16'd6788: out <= 16'hFFBA;    16'd6789: out <= 16'hFC65;    16'd6790: out <= 16'h0234;    16'd6791: out <= 16'h0BD8;
    16'd6792: out <= 16'h0425;    16'd6793: out <= 16'h00D9;    16'd6794: out <= 16'h05CB;    16'd6795: out <= 16'h0228;
    16'd6796: out <= 16'hFC65;    16'd6797: out <= 16'h0050;    16'd6798: out <= 16'h0BCE;    16'd6799: out <= 16'hFC32;
    16'd6800: out <= 16'h0335;    16'd6801: out <= 16'h03BD;    16'd6802: out <= 16'hFEFD;    16'd6803: out <= 16'h01E4;
    16'd6804: out <= 16'h027E;    16'd6805: out <= 16'h03D6;    16'd6806: out <= 16'h0162;    16'd6807: out <= 16'hF946;
    16'd6808: out <= 16'h062C;    16'd6809: out <= 16'h04A6;    16'd6810: out <= 16'h087E;    16'd6811: out <= 16'h05FE;
    16'd6812: out <= 16'h01C9;    16'd6813: out <= 16'h01F4;    16'd6814: out <= 16'h0359;    16'd6815: out <= 16'h027E;
    16'd6816: out <= 16'h024D;    16'd6817: out <= 16'h0783;    16'd6818: out <= 16'h036E;    16'd6819: out <= 16'h01D6;
    16'd6820: out <= 16'h0160;    16'd6821: out <= 16'h05CE;    16'd6822: out <= 16'h0061;    16'd6823: out <= 16'h0A67;
    16'd6824: out <= 16'h04A3;    16'd6825: out <= 16'hFCC9;    16'd6826: out <= 16'h010F;    16'd6827: out <= 16'hFFF6;
    16'd6828: out <= 16'h0507;    16'd6829: out <= 16'h07AB;    16'd6830: out <= 16'h0568;    16'd6831: out <= 16'h07D4;
    16'd6832: out <= 16'h0137;    16'd6833: out <= 16'h0399;    16'd6834: out <= 16'hFC84;    16'd6835: out <= 16'h07AC;
    16'd6836: out <= 16'h07EF;    16'd6837: out <= 16'h0330;    16'd6838: out <= 16'h06E8;    16'd6839: out <= 16'h003E;
    16'd6840: out <= 16'h07D4;    16'd6841: out <= 16'h005A;    16'd6842: out <= 16'h069A;    16'd6843: out <= 16'h08B0;
    16'd6844: out <= 16'h0256;    16'd6845: out <= 16'h049A;    16'd6846: out <= 16'h01EB;    16'd6847: out <= 16'h0661;
    16'd6848: out <= 16'h0AF5;    16'd6849: out <= 16'hFD5E;    16'd6850: out <= 16'h013D;    16'd6851: out <= 16'h090B;
    16'd6852: out <= 16'h02FE;    16'd6853: out <= 16'hFBD9;    16'd6854: out <= 16'hFCFB;    16'd6855: out <= 16'h001F;
    16'd6856: out <= 16'h04CC;    16'd6857: out <= 16'h032A;    16'd6858: out <= 16'h00B4;    16'd6859: out <= 16'h01B3;
    16'd6860: out <= 16'hFD8C;    16'd6861: out <= 16'h045E;    16'd6862: out <= 16'h0227;    16'd6863: out <= 16'h0873;
    16'd6864: out <= 16'hFD3C;    16'd6865: out <= 16'h04AE;    16'd6866: out <= 16'hFB68;    16'd6867: out <= 16'hFA27;
    16'd6868: out <= 16'hFDDF;    16'd6869: out <= 16'h06A5;    16'd6870: out <= 16'hFAD7;    16'd6871: out <= 16'h0636;
    16'd6872: out <= 16'h0551;    16'd6873: out <= 16'h052A;    16'd6874: out <= 16'hFBAB;    16'd6875: out <= 16'h0183;
    16'd6876: out <= 16'hFD39;    16'd6877: out <= 16'hF97A;    16'd6878: out <= 16'h00D8;    16'd6879: out <= 16'h01F6;
    16'd6880: out <= 16'hFDF0;    16'd6881: out <= 16'h04BD;    16'd6882: out <= 16'h01FC;    16'd6883: out <= 16'hF7E3;
    16'd6884: out <= 16'hFEF7;    16'd6885: out <= 16'hFBAC;    16'd6886: out <= 16'h07A0;    16'd6887: out <= 16'hFCB0;
    16'd6888: out <= 16'hFE07;    16'd6889: out <= 16'hFBE8;    16'd6890: out <= 16'hFA4E;    16'd6891: out <= 16'h001D;
    16'd6892: out <= 16'h0090;    16'd6893: out <= 16'h05B5;    16'd6894: out <= 16'h03E9;    16'd6895: out <= 16'h0730;
    16'd6896: out <= 16'hFA16;    16'd6897: out <= 16'hFE81;    16'd6898: out <= 16'hFFC4;    16'd6899: out <= 16'hFB33;
    16'd6900: out <= 16'h0175;    16'd6901: out <= 16'h022A;    16'd6902: out <= 16'hFFFA;    16'd6903: out <= 16'h0511;
    16'd6904: out <= 16'h0486;    16'd6905: out <= 16'h0145;    16'd6906: out <= 16'hFBEB;    16'd6907: out <= 16'hFE00;
    16'd6908: out <= 16'h05D3;    16'd6909: out <= 16'hFAAB;    16'd6910: out <= 16'h0463;    16'd6911: out <= 16'h0366;
    16'd6912: out <= 16'h07E8;    16'd6913: out <= 16'hFB7E;    16'd6914: out <= 16'hFD94;    16'd6915: out <= 16'hFF23;
    16'd6916: out <= 16'hFEDE;    16'd6917: out <= 16'h004C;    16'd6918: out <= 16'hF80E;    16'd6919: out <= 16'h016A;
    16'd6920: out <= 16'h0652;    16'd6921: out <= 16'h0AA2;    16'd6922: out <= 16'hFD20;    16'd6923: out <= 16'h0363;
    16'd6924: out <= 16'hFC56;    16'd6925: out <= 16'hFCCC;    16'd6926: out <= 16'hFB85;    16'd6927: out <= 16'hFFFA;
    16'd6928: out <= 16'h027D;    16'd6929: out <= 16'h005D;    16'd6930: out <= 16'hFE07;    16'd6931: out <= 16'hF8C2;
    16'd6932: out <= 16'hFDA6;    16'd6933: out <= 16'hFBBD;    16'd6934: out <= 16'h04A6;    16'd6935: out <= 16'h0168;
    16'd6936: out <= 16'h0368;    16'd6937: out <= 16'h0756;    16'd6938: out <= 16'hF68A;    16'd6939: out <= 16'h07D4;
    16'd6940: out <= 16'h02AD;    16'd6941: out <= 16'hFF26;    16'd6942: out <= 16'hFFA0;    16'd6943: out <= 16'hF9D4;
    16'd6944: out <= 16'h05FC;    16'd6945: out <= 16'h03B1;    16'd6946: out <= 16'hFDBA;    16'd6947: out <= 16'h00EF;
    16'd6948: out <= 16'h0391;    16'd6949: out <= 16'hFE92;    16'd6950: out <= 16'hFFB0;    16'd6951: out <= 16'hFDAC;
    16'd6952: out <= 16'hF488;    16'd6953: out <= 16'h025E;    16'd6954: out <= 16'h02F1;    16'd6955: out <= 16'hFC9A;
    16'd6956: out <= 16'h021B;    16'd6957: out <= 16'hFCFC;    16'd6958: out <= 16'h0115;    16'd6959: out <= 16'h009D;
    16'd6960: out <= 16'h04CE;    16'd6961: out <= 16'hFD3B;    16'd6962: out <= 16'h0781;    16'd6963: out <= 16'hFEE1;
    16'd6964: out <= 16'h06A4;    16'd6965: out <= 16'h06CC;    16'd6966: out <= 16'h062A;    16'd6967: out <= 16'h0622;
    16'd6968: out <= 16'h0BE1;    16'd6969: out <= 16'h0C47;    16'd6970: out <= 16'h00A9;    16'd6971: out <= 16'hFDA4;
    16'd6972: out <= 16'h049C;    16'd6973: out <= 16'h052A;    16'd6974: out <= 16'h061A;    16'd6975: out <= 16'h034E;
    16'd6976: out <= 16'h0411;    16'd6977: out <= 16'h0435;    16'd6978: out <= 16'h05B6;    16'd6979: out <= 16'hFDF5;
    16'd6980: out <= 16'h030F;    16'd6981: out <= 16'h04AE;    16'd6982: out <= 16'h0846;    16'd6983: out <= 16'h06A1;
    16'd6984: out <= 16'hFB74;    16'd6985: out <= 16'h01DB;    16'd6986: out <= 16'h0D06;    16'd6987: out <= 16'hFE35;
    16'd6988: out <= 16'h05E7;    16'd6989: out <= 16'hF836;    16'd6990: out <= 16'h0443;    16'd6991: out <= 16'h057B;
    16'd6992: out <= 16'h0577;    16'd6993: out <= 16'hFEE2;    16'd6994: out <= 16'h0150;    16'd6995: out <= 16'h00D7;
    16'd6996: out <= 16'h03D5;    16'd6997: out <= 16'hFE5B;    16'd6998: out <= 16'h0550;    16'd6999: out <= 16'hFED7;
    16'd7000: out <= 16'hFEF4;    16'd7001: out <= 16'h03C9;    16'd7002: out <= 16'h0B55;    16'd7003: out <= 16'h090A;
    16'd7004: out <= 16'h026B;    16'd7005: out <= 16'h04E3;    16'd7006: out <= 16'h0259;    16'd7007: out <= 16'h06BF;
    16'd7008: out <= 16'h0398;    16'd7009: out <= 16'h0303;    16'd7010: out <= 16'h0336;    16'd7011: out <= 16'h0457;
    16'd7012: out <= 16'h0395;    16'd7013: out <= 16'h0065;    16'd7014: out <= 16'hFF7B;    16'd7015: out <= 16'h0954;
    16'd7016: out <= 16'h0623;    16'd7017: out <= 16'h083C;    16'd7018: out <= 16'h0299;    16'd7019: out <= 16'h04F2;
    16'd7020: out <= 16'h0836;    16'd7021: out <= 16'h02E7;    16'd7022: out <= 16'hFFD4;    16'd7023: out <= 16'h0A80;
    16'd7024: out <= 16'h0388;    16'd7025: out <= 16'hFEA3;    16'd7026: out <= 16'h015D;    16'd7027: out <= 16'h07D3;
    16'd7028: out <= 16'h0820;    16'd7029: out <= 16'h008B;    16'd7030: out <= 16'h0657;    16'd7031: out <= 16'h07A9;
    16'd7032: out <= 16'hFFE2;    16'd7033: out <= 16'h0BA7;    16'd7034: out <= 16'h0C68;    16'd7035: out <= 16'h05AD;
    16'd7036: out <= 16'hFD7D;    16'd7037: out <= 16'h04B1;    16'd7038: out <= 16'h06D5;    16'd7039: out <= 16'h0096;
    16'd7040: out <= 16'h07B9;    16'd7041: out <= 16'h005F;    16'd7042: out <= 16'h04D4;    16'd7043: out <= 16'h06D2;
    16'd7044: out <= 16'h0704;    16'd7045: out <= 16'h04AF;    16'd7046: out <= 16'h0663;    16'd7047: out <= 16'h0ABC;
    16'd7048: out <= 16'h01E4;    16'd7049: out <= 16'hFF68;    16'd7050: out <= 16'h00A0;    16'd7051: out <= 16'h05C1;
    16'd7052: out <= 16'hFDFF;    16'd7053: out <= 16'h084B;    16'd7054: out <= 16'h091E;    16'd7055: out <= 16'h0128;
    16'd7056: out <= 16'h038B;    16'd7057: out <= 16'h04BA;    16'd7058: out <= 16'h0328;    16'd7059: out <= 16'h0474;
    16'd7060: out <= 16'h06EC;    16'd7061: out <= 16'h01FC;    16'd7062: out <= 16'h025D;    16'd7063: out <= 16'h0813;
    16'd7064: out <= 16'h01AD;    16'd7065: out <= 16'hFD97;    16'd7066: out <= 16'hFF61;    16'd7067: out <= 16'h02F5;
    16'd7068: out <= 16'h05E0;    16'd7069: out <= 16'h03DA;    16'd7070: out <= 16'hFF90;    16'd7071: out <= 16'h08DA;
    16'd7072: out <= 16'hFFBF;    16'd7073: out <= 16'h03EA;    16'd7074: out <= 16'h037F;    16'd7075: out <= 16'h00F5;
    16'd7076: out <= 16'hFD68;    16'd7077: out <= 16'h067A;    16'd7078: out <= 16'h0B31;    16'd7079: out <= 16'h04D5;
    16'd7080: out <= 16'h050A;    16'd7081: out <= 16'h080A;    16'd7082: out <= 16'h040B;    16'd7083: out <= 16'h026D;
    16'd7084: out <= 16'h0456;    16'd7085: out <= 16'h06B1;    16'd7086: out <= 16'hFFF5;    16'd7087: out <= 16'h0423;
    16'd7088: out <= 16'h016B;    16'd7089: out <= 16'hFE8F;    16'd7090: out <= 16'h0797;    16'd7091: out <= 16'h06CD;
    16'd7092: out <= 16'h0729;    16'd7093: out <= 16'h037A;    16'd7094: out <= 16'hFF14;    16'd7095: out <= 16'h0EDE;
    16'd7096: out <= 16'h06C8;    16'd7097: out <= 16'h08C6;    16'd7098: out <= 16'h057C;    16'd7099: out <= 16'h0156;
    16'd7100: out <= 16'h067B;    16'd7101: out <= 16'h0477;    16'd7102: out <= 16'h0969;    16'd7103: out <= 16'h0382;
    16'd7104: out <= 16'h0723;    16'd7105: out <= 16'h03E3;    16'd7106: out <= 16'h084D;    16'd7107: out <= 16'h06F1;
    16'd7108: out <= 16'h0790;    16'd7109: out <= 16'hFD7F;    16'd7110: out <= 16'h0138;    16'd7111: out <= 16'hFF4E;
    16'd7112: out <= 16'hF8FF;    16'd7113: out <= 16'h0495;    16'd7114: out <= 16'hFE60;    16'd7115: out <= 16'h031B;
    16'd7116: out <= 16'hFEE0;    16'd7117: out <= 16'h0195;    16'd7118: out <= 16'h01DF;    16'd7119: out <= 16'hFC3D;
    16'd7120: out <= 16'h022E;    16'd7121: out <= 16'h0173;    16'd7122: out <= 16'hFDA9;    16'd7123: out <= 16'h00DB;
    16'd7124: out <= 16'hFCF7;    16'd7125: out <= 16'h000D;    16'd7126: out <= 16'hFF73;    16'd7127: out <= 16'hFE3B;
    16'd7128: out <= 16'hFCC6;    16'd7129: out <= 16'hFF27;    16'd7130: out <= 16'hFEFB;    16'd7131: out <= 16'hFC46;
    16'd7132: out <= 16'h07A9;    16'd7133: out <= 16'h0146;    16'd7134: out <= 16'hF97C;    16'd7135: out <= 16'h025A;
    16'd7136: out <= 16'hFE41;    16'd7137: out <= 16'hFC3E;    16'd7138: out <= 16'h0036;    16'd7139: out <= 16'h0153;
    16'd7140: out <= 16'h0023;    16'd7141: out <= 16'h02F3;    16'd7142: out <= 16'h01C6;    16'd7143: out <= 16'h0305;
    16'd7144: out <= 16'h03A5;    16'd7145: out <= 16'hFE3E;    16'd7146: out <= 16'h0571;    16'd7147: out <= 16'h04E8;
    16'd7148: out <= 16'hFFC3;    16'd7149: out <= 16'hFC5A;    16'd7150: out <= 16'h003E;    16'd7151: out <= 16'h02B0;
    16'd7152: out <= 16'hFF46;    16'd7153: out <= 16'h0422;    16'd7154: out <= 16'hFF94;    16'd7155: out <= 16'hF7C3;
    16'd7156: out <= 16'h0213;    16'd7157: out <= 16'h00BA;    16'd7158: out <= 16'h017A;    16'd7159: out <= 16'hFDC8;
    16'd7160: out <= 16'h0395;    16'd7161: out <= 16'h0452;    16'd7162: out <= 16'hFC9B;    16'd7163: out <= 16'hFABB;
    16'd7164: out <= 16'hFA24;    16'd7165: out <= 16'h0050;    16'd7166: out <= 16'hFF27;    16'd7167: out <= 16'h020B;
    16'd7168: out <= 16'h0033;    16'd7169: out <= 16'h0BAB;    16'd7170: out <= 16'h081F;    16'd7171: out <= 16'hFA25;
    16'd7172: out <= 16'h024A;    16'd7173: out <= 16'hFB0E;    16'd7174: out <= 16'h0192;    16'd7175: out <= 16'h09AA;
    16'd7176: out <= 16'hFDED;    16'd7177: out <= 16'hFC66;    16'd7178: out <= 16'h03E9;    16'd7179: out <= 16'h03CC;
    16'd7180: out <= 16'h0045;    16'd7181: out <= 16'h0370;    16'd7182: out <= 16'hFAFD;    16'd7183: out <= 16'hFDD6;
    16'd7184: out <= 16'h02DB;    16'd7185: out <= 16'h0B18;    16'd7186: out <= 16'hFED2;    16'd7187: out <= 16'h048D;
    16'd7188: out <= 16'hFACF;    16'd7189: out <= 16'hFE0C;    16'd7190: out <= 16'h0451;    16'd7191: out <= 16'hFEE3;
    16'd7192: out <= 16'hFFF8;    16'd7193: out <= 16'hFF35;    16'd7194: out <= 16'h01D7;    16'd7195: out <= 16'h06E7;
    16'd7196: out <= 16'h006A;    16'd7197: out <= 16'h006D;    16'd7198: out <= 16'h05D1;    16'd7199: out <= 16'hFF1B;
    16'd7200: out <= 16'hFD34;    16'd7201: out <= 16'h0299;    16'd7202: out <= 16'hFAA0;    16'd7203: out <= 16'h0430;
    16'd7204: out <= 16'hFF9E;    16'd7205: out <= 16'h0226;    16'd7206: out <= 16'hFAB2;    16'd7207: out <= 16'h04B1;
    16'd7208: out <= 16'hFE08;    16'd7209: out <= 16'h0B54;    16'd7210: out <= 16'h0022;    16'd7211: out <= 16'h0581;
    16'd7212: out <= 16'hFC69;    16'd7213: out <= 16'hFF0F;    16'd7214: out <= 16'h03B0;    16'd7215: out <= 16'h0605;
    16'd7216: out <= 16'hFE89;    16'd7217: out <= 16'hFEF7;    16'd7218: out <= 16'h0434;    16'd7219: out <= 16'h01E4;
    16'd7220: out <= 16'hFC92;    16'd7221: out <= 16'h075D;    16'd7222: out <= 16'h05FE;    16'd7223: out <= 16'h041C;
    16'd7224: out <= 16'h02DC;    16'd7225: out <= 16'hFFE9;    16'd7226: out <= 16'h0547;    16'd7227: out <= 16'h01BF;
    16'd7228: out <= 16'h0653;    16'd7229: out <= 16'h04E3;    16'd7230: out <= 16'h029F;    16'd7231: out <= 16'h0840;
    16'd7232: out <= 16'hFCB3;    16'd7233: out <= 16'hFD47;    16'd7234: out <= 16'h01CB;    16'd7235: out <= 16'h0624;
    16'd7236: out <= 16'h0236;    16'd7237: out <= 16'h0135;    16'd7238: out <= 16'h0073;    16'd7239: out <= 16'h02D7;
    16'd7240: out <= 16'h07A9;    16'd7241: out <= 16'h077D;    16'd7242: out <= 16'h0E37;    16'd7243: out <= 16'h0751;
    16'd7244: out <= 16'h03FD;    16'd7245: out <= 16'h01CB;    16'd7246: out <= 16'h0957;    16'd7247: out <= 16'h0A23;
    16'd7248: out <= 16'h04FB;    16'd7249: out <= 16'h01A2;    16'd7250: out <= 16'hFEC3;    16'd7251: out <= 16'hFE16;
    16'd7252: out <= 16'hFFD7;    16'd7253: out <= 16'h083B;    16'd7254: out <= 16'h043C;    16'd7255: out <= 16'h03E6;
    16'd7256: out <= 16'h07B6;    16'd7257: out <= 16'h0883;    16'd7258: out <= 16'h0271;    16'd7259: out <= 16'h0A88;
    16'd7260: out <= 16'h056D;    16'd7261: out <= 16'h0032;    16'd7262: out <= 16'hFECF;    16'd7263: out <= 16'h0E30;
    16'd7264: out <= 16'h0EAF;    16'd7265: out <= 16'h055B;    16'd7266: out <= 16'h00B8;    16'd7267: out <= 16'h0445;
    16'd7268: out <= 16'h0475;    16'd7269: out <= 16'h07C7;    16'd7270: out <= 16'h01BE;    16'd7271: out <= 16'h0180;
    16'd7272: out <= 16'hFD51;    16'd7273: out <= 16'h0085;    16'd7274: out <= 16'h0999;    16'd7275: out <= 16'h04B7;
    16'd7276: out <= 16'h08F6;    16'd7277: out <= 16'h07D1;    16'd7278: out <= 16'h04A3;    16'd7279: out <= 16'hFF32;
    16'd7280: out <= 16'h0393;    16'd7281: out <= 16'h0796;    16'd7282: out <= 16'h06D0;    16'd7283: out <= 16'h027B;
    16'd7284: out <= 16'h0608;    16'd7285: out <= 16'h03C2;    16'd7286: out <= 16'hFDB9;    16'd7287: out <= 16'h0612;
    16'd7288: out <= 16'h0C30;    16'd7289: out <= 16'h02EA;    16'd7290: out <= 16'h0705;    16'd7291: out <= 16'h0497;
    16'd7292: out <= 16'h04B4;    16'd7293: out <= 16'h003B;    16'd7294: out <= 16'h080A;    16'd7295: out <= 16'h0A1D;
    16'd7296: out <= 16'h03B3;    16'd7297: out <= 16'h0C75;    16'd7298: out <= 16'h0540;    16'd7299: out <= 16'hFE8B;
    16'd7300: out <= 16'hFFAF;    16'd7301: out <= 16'h05C7;    16'd7302: out <= 16'h0B58;    16'd7303: out <= 16'h05A5;
    16'd7304: out <= 16'h01B5;    16'd7305: out <= 16'h04E6;    16'd7306: out <= 16'hFE0B;    16'd7307: out <= 16'h035F;
    16'd7308: out <= 16'h0710;    16'd7309: out <= 16'h0566;    16'd7310: out <= 16'h04E0;    16'd7311: out <= 16'h029F;
    16'd7312: out <= 16'h0058;    16'd7313: out <= 16'h030B;    16'd7314: out <= 16'hFF95;    16'd7315: out <= 16'h02FD;
    16'd7316: out <= 16'h00B8;    16'd7317: out <= 16'h03B8;    16'd7318: out <= 16'hFED0;    16'd7319: out <= 16'hFE65;
    16'd7320: out <= 16'h0015;    16'd7321: out <= 16'h04AE;    16'd7322: out <= 16'h052C;    16'd7323: out <= 16'h0011;
    16'd7324: out <= 16'h01C9;    16'd7325: out <= 16'h0B6D;    16'd7326: out <= 16'hFEC5;    16'd7327: out <= 16'h0357;
    16'd7328: out <= 16'h0029;    16'd7329: out <= 16'h0325;    16'd7330: out <= 16'h02F0;    16'd7331: out <= 16'h05E0;
    16'd7332: out <= 16'h0951;    16'd7333: out <= 16'h05A2;    16'd7334: out <= 16'h00F1;    16'd7335: out <= 16'h04FE;
    16'd7336: out <= 16'h08DE;    16'd7337: out <= 16'h074A;    16'd7338: out <= 16'h0BE1;    16'd7339: out <= 16'h05C9;
    16'd7340: out <= 16'h0444;    16'd7341: out <= 16'h07C5;    16'd7342: out <= 16'h03F7;    16'd7343: out <= 16'h025E;
    16'd7344: out <= 16'h0667;    16'd7345: out <= 16'h0C56;    16'd7346: out <= 16'h019B;    16'd7347: out <= 16'h03AF;
    16'd7348: out <= 16'h06ED;    16'd7349: out <= 16'hFCE3;    16'd7350: out <= 16'h0407;    16'd7351: out <= 16'h0268;
    16'd7352: out <= 16'h026A;    16'd7353: out <= 16'hFE76;    16'd7354: out <= 16'h041F;    16'd7355: out <= 16'h0A3B;
    16'd7356: out <= 16'hFD8D;    16'd7357: out <= 16'h059A;    16'd7358: out <= 16'h0165;    16'd7359: out <= 16'h00E2;
    16'd7360: out <= 16'hFBBF;    16'd7361: out <= 16'h0427;    16'd7362: out <= 16'h031D;    16'd7363: out <= 16'h00A6;
    16'd7364: out <= 16'h0294;    16'd7365: out <= 16'h056E;    16'd7366: out <= 16'h0408;    16'd7367: out <= 16'hF945;
    16'd7368: out <= 16'hFCCD;    16'd7369: out <= 16'hFE18;    16'd7370: out <= 16'hFF46;    16'd7371: out <= 16'hFBF3;
    16'd7372: out <= 16'h042E;    16'd7373: out <= 16'hFE52;    16'd7374: out <= 16'hFB72;    16'd7375: out <= 16'h02D9;
    16'd7376: out <= 16'h0193;    16'd7377: out <= 16'hFF4E;    16'd7378: out <= 16'h0684;    16'd7379: out <= 16'hFE0A;
    16'd7380: out <= 16'hFF05;    16'd7381: out <= 16'h02E3;    16'd7382: out <= 16'hFADF;    16'd7383: out <= 16'h011E;
    16'd7384: out <= 16'h0174;    16'd7385: out <= 16'h0152;    16'd7386: out <= 16'h06C5;    16'd7387: out <= 16'hF8BB;
    16'd7388: out <= 16'hF58B;    16'd7389: out <= 16'hFDE3;    16'd7390: out <= 16'h07E6;    16'd7391: out <= 16'h0445;
    16'd7392: out <= 16'hFE9C;    16'd7393: out <= 16'hFBBC;    16'd7394: out <= 16'h012C;    16'd7395: out <= 16'hFFBA;
    16'd7396: out <= 16'hFBD4;    16'd7397: out <= 16'hFC08;    16'd7398: out <= 16'hFC8F;    16'd7399: out <= 16'hFF97;
    16'd7400: out <= 16'h01B0;    16'd7401: out <= 16'hF63F;    16'd7402: out <= 16'hFA81;    16'd7403: out <= 16'h00C5;
    16'd7404: out <= 16'h0590;    16'd7405: out <= 16'h05B7;    16'd7406: out <= 16'h0218;    16'd7407: out <= 16'h03E1;
    16'd7408: out <= 16'hFDCE;    16'd7409: out <= 16'h0A95;    16'd7410: out <= 16'h01F6;    16'd7411: out <= 16'hFAF8;
    16'd7412: out <= 16'h0116;    16'd7413: out <= 16'hFB08;    16'd7414: out <= 16'h0205;    16'd7415: out <= 16'h03AC;
    16'd7416: out <= 16'hFEA7;    16'd7417: out <= 16'h0869;    16'd7418: out <= 16'h073D;    16'd7419: out <= 16'h0403;
    16'd7420: out <= 16'h00DF;    16'd7421: out <= 16'h027B;    16'd7422: out <= 16'h0502;    16'd7423: out <= 16'h0101;
    16'd7424: out <= 16'hFFE3;    16'd7425: out <= 16'hFF61;    16'd7426: out <= 16'h0190;    16'd7427: out <= 16'hFF37;
    16'd7428: out <= 16'hFDA5;    16'd7429: out <= 16'hFF98;    16'd7430: out <= 16'h05DA;    16'd7431: out <= 16'h00F8;
    16'd7432: out <= 16'hFE36;    16'd7433: out <= 16'h0542;    16'd7434: out <= 16'hFD75;    16'd7435: out <= 16'h0241;
    16'd7436: out <= 16'hFC94;    16'd7437: out <= 16'h00EA;    16'd7438: out <= 16'hFEA5;    16'd7439: out <= 16'h013C;
    16'd7440: out <= 16'hFEB0;    16'd7441: out <= 16'h07E2;    16'd7442: out <= 16'hFA9E;    16'd7443: out <= 16'h04AA;
    16'd7444: out <= 16'hF61D;    16'd7445: out <= 16'h01EA;    16'd7446: out <= 16'h03C6;    16'd7447: out <= 16'hFF5D;
    16'd7448: out <= 16'h02EA;    16'd7449: out <= 16'hFD1C;    16'd7450: out <= 16'hFC8D;    16'd7451: out <= 16'h0261;
    16'd7452: out <= 16'h0235;    16'd7453: out <= 16'hFAEB;    16'd7454: out <= 16'h04FE;    16'd7455: out <= 16'hFFD2;
    16'd7456: out <= 16'h06D6;    16'd7457: out <= 16'hFF90;    16'd7458: out <= 16'h0911;    16'd7459: out <= 16'h0596;
    16'd7460: out <= 16'hFEC3;    16'd7461: out <= 16'h011A;    16'd7462: out <= 16'h00C3;    16'd7463: out <= 16'hFC8F;
    16'd7464: out <= 16'hFFEA;    16'd7465: out <= 16'h038B;    16'd7466: out <= 16'hFBE9;    16'd7467: out <= 16'h0786;
    16'd7468: out <= 16'hF9DC;    16'd7469: out <= 16'h063C;    16'd7470: out <= 16'h004F;    16'd7471: out <= 16'hFF3B;
    16'd7472: out <= 16'h0387;    16'd7473: out <= 16'hF9AA;    16'd7474: out <= 16'h03B2;    16'd7475: out <= 16'h01A6;
    16'd7476: out <= 16'h069C;    16'd7477: out <= 16'hFE9B;    16'd7478: out <= 16'h08A5;    16'd7479: out <= 16'h0456;
    16'd7480: out <= 16'h0772;    16'd7481: out <= 16'hFE91;    16'd7482: out <= 16'h0280;    16'd7483: out <= 16'h09FC;
    16'd7484: out <= 16'h02A2;    16'd7485: out <= 16'h04D2;    16'd7486: out <= 16'h0614;    16'd7487: out <= 16'h0458;
    16'd7488: out <= 16'h01DF;    16'd7489: out <= 16'h03BA;    16'd7490: out <= 16'h0406;    16'd7491: out <= 16'h01A9;
    16'd7492: out <= 16'hFDAA;    16'd7493: out <= 16'h07D8;    16'd7494: out <= 16'h05DF;    16'd7495: out <= 16'h0185;
    16'd7496: out <= 16'hFFBE;    16'd7497: out <= 16'hFDE5;    16'd7498: out <= 16'h05A5;    16'd7499: out <= 16'h0421;
    16'd7500: out <= 16'hFFC6;    16'd7501: out <= 16'h08A0;    16'd7502: out <= 16'h0479;    16'd7503: out <= 16'h042D;
    16'd7504: out <= 16'h0638;    16'd7505: out <= 16'h0359;    16'd7506: out <= 16'h00D3;    16'd7507: out <= 16'hFCF3;
    16'd7508: out <= 16'h0237;    16'd7509: out <= 16'h0562;    16'd7510: out <= 16'h0600;    16'd7511: out <= 16'h04EA;
    16'd7512: out <= 16'h0240;    16'd7513: out <= 16'h08E7;    16'd7514: out <= 16'hFB7E;    16'd7515: out <= 16'h01A1;
    16'd7516: out <= 16'h08CD;    16'd7517: out <= 16'h0A36;    16'd7518: out <= 16'h00AA;    16'd7519: out <= 16'h04A6;
    16'd7520: out <= 16'h028D;    16'd7521: out <= 16'h0677;    16'd7522: out <= 16'h085F;    16'd7523: out <= 16'hFFA7;
    16'd7524: out <= 16'h0297;    16'd7525: out <= 16'h0041;    16'd7526: out <= 16'h04AB;    16'd7527: out <= 16'h007B;
    16'd7528: out <= 16'h04EB;    16'd7529: out <= 16'h022F;    16'd7530: out <= 16'h0637;    16'd7531: out <= 16'h0805;
    16'd7532: out <= 16'h0237;    16'd7533: out <= 16'h0435;    16'd7534: out <= 16'h06C4;    16'd7535: out <= 16'h00D4;
    16'd7536: out <= 16'h0346;    16'd7537: out <= 16'h0815;    16'd7538: out <= 16'h01C1;    16'd7539: out <= 16'hFAFD;
    16'd7540: out <= 16'h014A;    16'd7541: out <= 16'h015A;    16'd7542: out <= 16'h05CA;    16'd7543: out <= 16'h0181;
    16'd7544: out <= 16'h079B;    16'd7545: out <= 16'h06F3;    16'd7546: out <= 16'h047E;    16'd7547: out <= 16'h02DC;
    16'd7548: out <= 16'h062C;    16'd7549: out <= 16'h0602;    16'd7550: out <= 16'h00D5;    16'd7551: out <= 16'h0A69;
    16'd7552: out <= 16'h04AA;    16'd7553: out <= 16'h013E;    16'd7554: out <= 16'h076F;    16'd7555: out <= 16'h037F;
    16'd7556: out <= 16'h073B;    16'd7557: out <= 16'h067C;    16'd7558: out <= 16'hFF73;    16'd7559: out <= 16'h066D;
    16'd7560: out <= 16'h08CF;    16'd7561: out <= 16'h0061;    16'd7562: out <= 16'h0444;    16'd7563: out <= 16'h03CA;
    16'd7564: out <= 16'h0705;    16'd7565: out <= 16'h0453;    16'd7566: out <= 16'h0197;    16'd7567: out <= 16'hFFAC;
    16'd7568: out <= 16'h0332;    16'd7569: out <= 16'hFD8C;    16'd7570: out <= 16'h0771;    16'd7571: out <= 16'h052D;
    16'd7572: out <= 16'hFF7F;    16'd7573: out <= 16'h0807;    16'd7574: out <= 16'h0318;    16'd7575: out <= 16'h07AC;
    16'd7576: out <= 16'h04C7;    16'd7577: out <= 16'h051F;    16'd7578: out <= 16'h031C;    16'd7579: out <= 16'h0553;
    16'd7580: out <= 16'h083D;    16'd7581: out <= 16'h0599;    16'd7582: out <= 16'h0389;    16'd7583: out <= 16'h00F9;
    16'd7584: out <= 16'h0083;    16'd7585: out <= 16'h07A7;    16'd7586: out <= 16'h05C3;    16'd7587: out <= 16'h0715;
    16'd7588: out <= 16'h08F1;    16'd7589: out <= 16'h0569;    16'd7590: out <= 16'h04E2;    16'd7591: out <= 16'hFD24;
    16'd7592: out <= 16'hFED4;    16'd7593: out <= 16'hFED3;    16'd7594: out <= 16'h0194;    16'd7595: out <= 16'h0753;
    16'd7596: out <= 16'h051F;    16'd7597: out <= 16'h0A1C;    16'd7598: out <= 16'h092D;    16'd7599: out <= 16'h070F;
    16'd7600: out <= 16'h03BB;    16'd7601: out <= 16'h0221;    16'd7602: out <= 16'h0479;    16'd7603: out <= 16'h02E5;
    16'd7604: out <= 16'h00BE;    16'd7605: out <= 16'h01BD;    16'd7606: out <= 16'h0175;    16'd7607: out <= 16'h0025;
    16'd7608: out <= 16'hFFE4;    16'd7609: out <= 16'h06D4;    16'd7610: out <= 16'h0720;    16'd7611: out <= 16'hFD00;
    16'd7612: out <= 16'hFDD6;    16'd7613: out <= 16'h0B00;    16'd7614: out <= 16'h08C5;    16'd7615: out <= 16'h049E;
    16'd7616: out <= 16'h0848;    16'd7617: out <= 16'h0848;    16'd7618: out <= 16'hFA17;    16'd7619: out <= 16'h0554;
    16'd7620: out <= 16'h03FE;    16'd7621: out <= 16'h0134;    16'd7622: out <= 16'h02F2;    16'd7623: out <= 16'hFF18;
    16'd7624: out <= 16'h0389;    16'd7625: out <= 16'h0099;    16'd7626: out <= 16'h0522;    16'd7627: out <= 16'h03A9;
    16'd7628: out <= 16'h0034;    16'd7629: out <= 16'h04AD;    16'd7630: out <= 16'hFB53;    16'd7631: out <= 16'h01E1;
    16'd7632: out <= 16'h0084;    16'd7633: out <= 16'hF9AD;    16'd7634: out <= 16'hFFC1;    16'd7635: out <= 16'h0183;
    16'd7636: out <= 16'hFE1A;    16'd7637: out <= 16'h05C2;    16'd7638: out <= 16'hFF66;    16'd7639: out <= 16'h0054;
    16'd7640: out <= 16'h04F7;    16'd7641: out <= 16'hFEEF;    16'd7642: out <= 16'hFE7B;    16'd7643: out <= 16'hFA13;
    16'd7644: out <= 16'h02AC;    16'd7645: out <= 16'h00C7;    16'd7646: out <= 16'h0006;    16'd7647: out <= 16'h00AD;
    16'd7648: out <= 16'h002B;    16'd7649: out <= 16'h027C;    16'd7650: out <= 16'h06F5;    16'd7651: out <= 16'hFAEC;
    16'd7652: out <= 16'h05C2;    16'd7653: out <= 16'hFAC9;    16'd7654: out <= 16'hFEC1;    16'd7655: out <= 16'h03BB;
    16'd7656: out <= 16'h007D;    16'd7657: out <= 16'h064C;    16'd7658: out <= 16'h027F;    16'd7659: out <= 16'h0112;
    16'd7660: out <= 16'hFC56;    16'd7661: out <= 16'h034B;    16'd7662: out <= 16'hFED0;    16'd7663: out <= 16'h03F6;
    16'd7664: out <= 16'hFDA1;    16'd7665: out <= 16'hF5B4;    16'd7666: out <= 16'h02D7;    16'd7667: out <= 16'h0030;
    16'd7668: out <= 16'h044B;    16'd7669: out <= 16'h0467;    16'd7670: out <= 16'hF868;    16'd7671: out <= 16'h0188;
    16'd7672: out <= 16'hFF34;    16'd7673: out <= 16'hFF93;    16'd7674: out <= 16'hFF88;    16'd7675: out <= 16'hFB0C;
    16'd7676: out <= 16'h0217;    16'd7677: out <= 16'h0013;    16'd7678: out <= 16'h039D;    16'd7679: out <= 16'h02B4;
    16'd7680: out <= 16'hFDE0;    16'd7681: out <= 16'h03FB;    16'd7682: out <= 16'hFD46;    16'd7683: out <= 16'h0A2E;
    16'd7684: out <= 16'hFA91;    16'd7685: out <= 16'h00EB;    16'd7686: out <= 16'h0589;    16'd7687: out <= 16'h02DC;
    16'd7688: out <= 16'h029F;    16'd7689: out <= 16'h06B7;    16'd7690: out <= 16'hFDD8;    16'd7691: out <= 16'h0085;
    16'd7692: out <= 16'hFA35;    16'd7693: out <= 16'hFEA3;    16'd7694: out <= 16'h05C5;    16'd7695: out <= 16'h0324;
    16'd7696: out <= 16'hFC67;    16'd7697: out <= 16'h0250;    16'd7698: out <= 16'h05D0;    16'd7699: out <= 16'hFF7B;
    16'd7700: out <= 16'hFFE2;    16'd7701: out <= 16'h007C;    16'd7702: out <= 16'hFB2A;    16'd7703: out <= 16'hF8F8;
    16'd7704: out <= 16'h012E;    16'd7705: out <= 16'h00C4;    16'd7706: out <= 16'h0017;    16'd7707: out <= 16'hFFB8;
    16'd7708: out <= 16'hFE1A;    16'd7709: out <= 16'h04F5;    16'd7710: out <= 16'h04BE;    16'd7711: out <= 16'h03FD;
    16'd7712: out <= 16'hFAA9;    16'd7713: out <= 16'h0346;    16'd7714: out <= 16'hFFF7;    16'd7715: out <= 16'hFF34;
    16'd7716: out <= 16'h0334;    16'd7717: out <= 16'hFED4;    16'd7718: out <= 16'h03BF;    16'd7719: out <= 16'hFE66;
    16'd7720: out <= 16'hFB96;    16'd7721: out <= 16'hFE2B;    16'd7722: out <= 16'h08C5;    16'd7723: out <= 16'h0178;
    16'd7724: out <= 16'h0458;    16'd7725: out <= 16'h05F5;    16'd7726: out <= 16'hFC91;    16'd7727: out <= 16'hFA56;
    16'd7728: out <= 16'h0278;    16'd7729: out <= 16'hFF70;    16'd7730: out <= 16'h01D7;    16'd7731: out <= 16'hFE2C;
    16'd7732: out <= 16'h0458;    16'd7733: out <= 16'h03B1;    16'd7734: out <= 16'h035E;    16'd7735: out <= 16'h043E;
    16'd7736: out <= 16'h025B;    16'd7737: out <= 16'h001C;    16'd7738: out <= 16'hFD32;    16'd7739: out <= 16'h0322;
    16'd7740: out <= 16'h00C0;    16'd7741: out <= 16'h0A33;    16'd7742: out <= 16'h086F;    16'd7743: out <= 16'h007D;
    16'd7744: out <= 16'h0121;    16'd7745: out <= 16'hFB8D;    16'd7746: out <= 16'h0964;    16'd7747: out <= 16'h07E8;
    16'd7748: out <= 16'hFE83;    16'd7749: out <= 16'h0A29;    16'd7750: out <= 16'h04DB;    16'd7751: out <= 16'h0526;
    16'd7752: out <= 16'h0683;    16'd7753: out <= 16'h0373;    16'd7754: out <= 16'h06A0;    16'd7755: out <= 16'h006A;
    16'd7756: out <= 16'hFF5E;    16'd7757: out <= 16'h0648;    16'd7758: out <= 16'h043D;    16'd7759: out <= 16'h04E4;
    16'd7760: out <= 16'hFFE8;    16'd7761: out <= 16'h0106;    16'd7762: out <= 16'h0705;    16'd7763: out <= 16'h05BD;
    16'd7764: out <= 16'h070D;    16'd7765: out <= 16'h0185;    16'd7766: out <= 16'hFFCE;    16'd7767: out <= 16'h0414;
    16'd7768: out <= 16'h0B3E;    16'd7769: out <= 16'h0823;    16'd7770: out <= 16'h051B;    16'd7771: out <= 16'hFFEE;
    16'd7772: out <= 16'h08D5;    16'd7773: out <= 16'h0358;    16'd7774: out <= 16'h0281;    16'd7775: out <= 16'hFCF0;
    16'd7776: out <= 16'hFE3C;    16'd7777: out <= 16'h0545;    16'd7778: out <= 16'hFF94;    16'd7779: out <= 16'hFB61;
    16'd7780: out <= 16'hFC9C;    16'd7781: out <= 16'h0023;    16'd7782: out <= 16'h0782;    16'd7783: out <= 16'hFDFF;
    16'd7784: out <= 16'h014A;    16'd7785: out <= 16'h043F;    16'd7786: out <= 16'h00B4;    16'd7787: out <= 16'h02C9;
    16'd7788: out <= 16'h0948;    16'd7789: out <= 16'h019C;    16'd7790: out <= 16'h0AC5;    16'd7791: out <= 16'h005B;
    16'd7792: out <= 16'h028F;    16'd7793: out <= 16'h08C5;    16'd7794: out <= 16'h0254;    16'd7795: out <= 16'h06BC;
    16'd7796: out <= 16'hFED8;    16'd7797: out <= 16'hFECF;    16'd7798: out <= 16'h01F3;    16'd7799: out <= 16'h047F;
    16'd7800: out <= 16'hFFAE;    16'd7801: out <= 16'h04F7;    16'd7802: out <= 16'h0090;    16'd7803: out <= 16'h0043;
    16'd7804: out <= 16'h03E5;    16'd7805: out <= 16'h07F7;    16'd7806: out <= 16'h04B6;    16'd7807: out <= 16'h0104;
    16'd7808: out <= 16'hFE70;    16'd7809: out <= 16'h033F;    16'd7810: out <= 16'h06E7;    16'd7811: out <= 16'h0B99;
    16'd7812: out <= 16'h042B;    16'd7813: out <= 16'h0544;    16'd7814: out <= 16'h032C;    16'd7815: out <= 16'hFF76;
    16'd7816: out <= 16'hFF9C;    16'd7817: out <= 16'h0645;    16'd7818: out <= 16'h02AE;    16'd7819: out <= 16'h0453;
    16'd7820: out <= 16'h00CF;    16'd7821: out <= 16'h0468;    16'd7822: out <= 16'h0790;    16'd7823: out <= 16'hFDAE;
    16'd7824: out <= 16'h00BC;    16'd7825: out <= 16'hFA17;    16'd7826: out <= 16'h0154;    16'd7827: out <= 16'hFF71;
    16'd7828: out <= 16'h037E;    16'd7829: out <= 16'h041C;    16'd7830: out <= 16'h06E4;    16'd7831: out <= 16'h054D;
    16'd7832: out <= 16'h06EF;    16'd7833: out <= 16'h01D4;    16'd7834: out <= 16'hFF50;    16'd7835: out <= 16'h08F7;
    16'd7836: out <= 16'hFD3C;    16'd7837: out <= 16'h0873;    16'd7838: out <= 16'h056C;    16'd7839: out <= 16'h07F6;
    16'd7840: out <= 16'h048F;    16'd7841: out <= 16'h06F6;    16'd7842: out <= 16'hFF39;    16'd7843: out <= 16'h0477;
    16'd7844: out <= 16'hFD78;    16'd7845: out <= 16'h036B;    16'd7846: out <= 16'h0A99;    16'd7847: out <= 16'hFFC7;
    16'd7848: out <= 16'h0AE0;    16'd7849: out <= 16'h06CE;    16'd7850: out <= 16'h053C;    16'd7851: out <= 16'h05E5;
    16'd7852: out <= 16'h06F7;    16'd7853: out <= 16'hFEFC;    16'd7854: out <= 16'hFE51;    16'd7855: out <= 16'h067E;
    16'd7856: out <= 16'h0175;    16'd7857: out <= 16'h0222;    16'd7858: out <= 16'h06E0;    16'd7859: out <= 16'h01EF;
    16'd7860: out <= 16'h027E;    16'd7861: out <= 16'hFC03;    16'd7862: out <= 16'h0275;    16'd7863: out <= 16'hFF4F;
    16'd7864: out <= 16'h01FF;    16'd7865: out <= 16'h018E;    16'd7866: out <= 16'h03AF;    16'd7867: out <= 16'h06B3;
    16'd7868: out <= 16'h04A3;    16'd7869: out <= 16'h0089;    16'd7870: out <= 16'h0A2B;    16'd7871: out <= 16'hFA33;
    16'd7872: out <= 16'hFACC;    16'd7873: out <= 16'h03DD;    16'd7874: out <= 16'h02C8;    16'd7875: out <= 16'hFCF9;
    16'd7876: out <= 16'h0B22;    16'd7877: out <= 16'h01FE;    16'd7878: out <= 16'h0451;    16'd7879: out <= 16'hFF60;
    16'd7880: out <= 16'h0458;    16'd7881: out <= 16'hFF1B;    16'd7882: out <= 16'h00E6;    16'd7883: out <= 16'h0105;
    16'd7884: out <= 16'h0244;    16'd7885: out <= 16'hFBC9;    16'd7886: out <= 16'h0256;    16'd7887: out <= 16'h02D0;
    16'd7888: out <= 16'hF9F1;    16'd7889: out <= 16'hFF7F;    16'd7890: out <= 16'h0232;    16'd7891: out <= 16'hFD81;
    16'd7892: out <= 16'hFBE1;    16'd7893: out <= 16'hFEBE;    16'd7894: out <= 16'hFAC6;    16'd7895: out <= 16'hFA73;
    16'd7896: out <= 16'hFE4F;    16'd7897: out <= 16'h0452;    16'd7898: out <= 16'h007C;    16'd7899: out <= 16'hFEC6;
    16'd7900: out <= 16'hFEC3;    16'd7901: out <= 16'hFAFA;    16'd7902: out <= 16'h0398;    16'd7903: out <= 16'h037E;
    16'd7904: out <= 16'hFB2A;    16'd7905: out <= 16'hFB2C;    16'd7906: out <= 16'h0155;    16'd7907: out <= 16'hFD4D;
    16'd7908: out <= 16'h0402;    16'd7909: out <= 16'hFFF4;    16'd7910: out <= 16'h00A2;    16'd7911: out <= 16'hFD78;
    16'd7912: out <= 16'h0345;    16'd7913: out <= 16'h0254;    16'd7914: out <= 16'h0236;    16'd7915: out <= 16'h025C;
    16'd7916: out <= 16'hFA89;    16'd7917: out <= 16'h00C7;    16'd7918: out <= 16'h01CB;    16'd7919: out <= 16'h0059;
    16'd7920: out <= 16'h01F6;    16'd7921: out <= 16'hFE8C;    16'd7922: out <= 16'hFE89;    16'd7923: out <= 16'h015E;
    16'd7924: out <= 16'hFEDF;    16'd7925: out <= 16'h028C;    16'd7926: out <= 16'h0089;    16'd7927: out <= 16'hFAD2;
    16'd7928: out <= 16'h061F;    16'd7929: out <= 16'hFC46;    16'd7930: out <= 16'h0002;    16'd7931: out <= 16'h02A5;
    16'd7932: out <= 16'hF878;    16'd7933: out <= 16'hFDF8;    16'd7934: out <= 16'hFE50;    16'd7935: out <= 16'hFDE0;
    16'd7936: out <= 16'hFFBA;    16'd7937: out <= 16'h02DE;    16'd7938: out <= 16'hF79F;    16'd7939: out <= 16'h002E;
    16'd7940: out <= 16'hFE60;    16'd7941: out <= 16'hFFF7;    16'd7942: out <= 16'h041C;    16'd7943: out <= 16'hFCEA;
    16'd7944: out <= 16'hFF42;    16'd7945: out <= 16'hFED7;    16'd7946: out <= 16'h0259;    16'd7947: out <= 16'hFA4E;
    16'd7948: out <= 16'hFC28;    16'd7949: out <= 16'hF9F2;    16'd7950: out <= 16'hFF76;    16'd7951: out <= 16'h02EA;
    16'd7952: out <= 16'h0246;    16'd7953: out <= 16'h0486;    16'd7954: out <= 16'h087C;    16'd7955: out <= 16'h0217;
    16'd7956: out <= 16'hFE50;    16'd7957: out <= 16'hFC81;    16'd7958: out <= 16'hFF88;    16'd7959: out <= 16'hFEC7;
    16'd7960: out <= 16'h06E8;    16'd7961: out <= 16'hFDE2;    16'd7962: out <= 16'h003A;    16'd7963: out <= 16'h048F;
    16'd7964: out <= 16'h01DF;    16'd7965: out <= 16'h0062;    16'd7966: out <= 16'hF912;    16'd7967: out <= 16'h00C4;
    16'd7968: out <= 16'hFE09;    16'd7969: out <= 16'hFB55;    16'd7970: out <= 16'h02D5;    16'd7971: out <= 16'hFC17;
    16'd7972: out <= 16'hFC2B;    16'd7973: out <= 16'hFACE;    16'd7974: out <= 16'hFEF3;    16'd7975: out <= 16'hFFA1;
    16'd7976: out <= 16'h026E;    16'd7977: out <= 16'h01F1;    16'd7978: out <= 16'h0066;    16'd7979: out <= 16'h019A;
    16'd7980: out <= 16'h01BB;    16'd7981: out <= 16'h0324;    16'd7982: out <= 16'hFCBB;    16'd7983: out <= 16'hFDFB;
    16'd7984: out <= 16'hFCC6;    16'd7985: out <= 16'h0727;    16'd7986: out <= 16'h0A7B;    16'd7987: out <= 16'h09F4;
    16'd7988: out <= 16'h03BF;    16'd7989: out <= 16'hFDE6;    16'd7990: out <= 16'h0065;    16'd7991: out <= 16'h068A;
    16'd7992: out <= 16'h09E5;    16'd7993: out <= 16'h0B1A;    16'd7994: out <= 16'h05B7;    16'd7995: out <= 16'h082B;
    16'd7996: out <= 16'h024E;    16'd7997: out <= 16'hFDE4;    16'd7998: out <= 16'h004E;    16'd7999: out <= 16'h057C;
    16'd8000: out <= 16'h03D4;    16'd8001: out <= 16'h006F;    16'd8002: out <= 16'h0728;    16'd8003: out <= 16'h007E;
    16'd8004: out <= 16'h05A5;    16'd8005: out <= 16'h05D0;    16'd8006: out <= 16'h09CA;    16'd8007: out <= 16'h0712;
    16'd8008: out <= 16'hFCC8;    16'd8009: out <= 16'h0748;    16'd8010: out <= 16'h04EC;    16'd8011: out <= 16'h0CEC;
    16'd8012: out <= 16'h04FB;    16'd8013: out <= 16'h04B7;    16'd8014: out <= 16'h02DD;    16'd8015: out <= 16'h09FF;
    16'd8016: out <= 16'hFD04;    16'd8017: out <= 16'h0451;    16'd8018: out <= 16'h0107;    16'd8019: out <= 16'h0215;
    16'd8020: out <= 16'h076A;    16'd8021: out <= 16'h05D2;    16'd8022: out <= 16'h0017;    16'd8023: out <= 16'h028F;
    16'd8024: out <= 16'hFDC6;    16'd8025: out <= 16'h0704;    16'd8026: out <= 16'h0814;    16'd8027: out <= 16'h0572;
    16'd8028: out <= 16'h003E;    16'd8029: out <= 16'h098D;    16'd8030: out <= 16'hFF9C;    16'd8031: out <= 16'h0837;
    16'd8032: out <= 16'h01AA;    16'd8033: out <= 16'h0F64;    16'd8034: out <= 16'h07E5;    16'd8035: out <= 16'h0303;
    16'd8036: out <= 16'h053B;    16'd8037: out <= 16'h04D2;    16'd8038: out <= 16'h03D5;    16'd8039: out <= 16'h01A7;
    16'd8040: out <= 16'h0686;    16'd8041: out <= 16'h01C5;    16'd8042: out <= 16'h0532;    16'd8043: out <= 16'h0396;
    16'd8044: out <= 16'h0341;    16'd8045: out <= 16'h005D;    16'd8046: out <= 16'h034F;    16'd8047: out <= 16'h04DC;
    16'd8048: out <= 16'h01E9;    16'd8049: out <= 16'hFB38;    16'd8050: out <= 16'h0750;    16'd8051: out <= 16'h0ABD;
    16'd8052: out <= 16'h0320;    16'd8053: out <= 16'h03C6;    16'd8054: out <= 16'h0527;    16'd8055: out <= 16'hFD2B;
    16'd8056: out <= 16'h03F3;    16'd8057: out <= 16'h00B4;    16'd8058: out <= 16'h0691;    16'd8059: out <= 16'h02C5;
    16'd8060: out <= 16'h0527;    16'd8061: out <= 16'h0238;    16'd8062: out <= 16'hFBEA;    16'd8063: out <= 16'hFE35;
    16'd8064: out <= 16'h02B8;    16'd8065: out <= 16'h0556;    16'd8066: out <= 16'h0190;    16'd8067: out <= 16'h0577;
    16'd8068: out <= 16'h059B;    16'd8069: out <= 16'h0422;    16'd8070: out <= 16'hFF9B;    16'd8071: out <= 16'h0480;
    16'd8072: out <= 16'h04C7;    16'd8073: out <= 16'h040D;    16'd8074: out <= 16'h0B83;    16'd8075: out <= 16'h0293;
    16'd8076: out <= 16'h02DF;    16'd8077: out <= 16'h062D;    16'd8078: out <= 16'h03A3;    16'd8079: out <= 16'h0628;
    16'd8080: out <= 16'h0739;    16'd8081: out <= 16'h04E1;    16'd8082: out <= 16'hFFA6;    16'd8083: out <= 16'h0686;
    16'd8084: out <= 16'hFEB8;    16'd8085: out <= 16'hFF51;    16'd8086: out <= 16'h0B48;    16'd8087: out <= 16'h0317;
    16'd8088: out <= 16'h07C0;    16'd8089: out <= 16'h0B07;    16'd8090: out <= 16'h05DE;    16'd8091: out <= 16'h0244;
    16'd8092: out <= 16'h03F1;    16'd8093: out <= 16'h023E;    16'd8094: out <= 16'h06AC;    16'd8095: out <= 16'h0253;
    16'd8096: out <= 16'hFFE6;    16'd8097: out <= 16'h0262;    16'd8098: out <= 16'h031F;    16'd8099: out <= 16'h0270;
    16'd8100: out <= 16'h0659;    16'd8101: out <= 16'h0102;    16'd8102: out <= 16'h01D3;    16'd8103: out <= 16'h08E7;
    16'd8104: out <= 16'h05FB;    16'd8105: out <= 16'h0160;    16'd8106: out <= 16'h092F;    16'd8107: out <= 16'h0001;
    16'd8108: out <= 16'h0387;    16'd8109: out <= 16'h0344;    16'd8110: out <= 16'h0C5F;    16'd8111: out <= 16'h015D;
    16'd8112: out <= 16'h0068;    16'd8113: out <= 16'h06D1;    16'd8114: out <= 16'h05F6;    16'd8115: out <= 16'hFEE9;
    16'd8116: out <= 16'hFE06;    16'd8117: out <= 16'h050F;    16'd8118: out <= 16'h034C;    16'd8119: out <= 16'h06E5;
    16'd8120: out <= 16'hFE3C;    16'd8121: out <= 16'h0143;    16'd8122: out <= 16'hFE70;    16'd8123: out <= 16'h027E;
    16'd8124: out <= 16'h0924;    16'd8125: out <= 16'h0777;    16'd8126: out <= 16'h041B;    16'd8127: out <= 16'h0460;
    16'd8128: out <= 16'h04A3;    16'd8129: out <= 16'h014F;    16'd8130: out <= 16'h04F0;    16'd8131: out <= 16'h063E;
    16'd8132: out <= 16'h059B;    16'd8133: out <= 16'h09E6;    16'd8134: out <= 16'h070E;    16'd8135: out <= 16'h02FE;
    16'd8136: out <= 16'h044D;    16'd8137: out <= 16'h0477;    16'd8138: out <= 16'h0196;    16'd8139: out <= 16'h039E;
    16'd8140: out <= 16'hFE17;    16'd8141: out <= 16'h0171;    16'd8142: out <= 16'hF9CC;    16'd8143: out <= 16'hFEE8;
    16'd8144: out <= 16'hFD48;    16'd8145: out <= 16'hFFB6;    16'd8146: out <= 16'hFD93;    16'd8147: out <= 16'hFBEE;
    16'd8148: out <= 16'h0284;    16'd8149: out <= 16'hF8A1;    16'd8150: out <= 16'h0204;    16'd8151: out <= 16'h03FC;
    16'd8152: out <= 16'hF8EF;    16'd8153: out <= 16'h02E3;    16'd8154: out <= 16'hFEC9;    16'd8155: out <= 16'h00EE;
    16'd8156: out <= 16'h02B3;    16'd8157: out <= 16'h02C5;    16'd8158: out <= 16'hFEC6;    16'd8159: out <= 16'hFFD0;
    16'd8160: out <= 16'hF89F;    16'd8161: out <= 16'hFC55;    16'd8162: out <= 16'hFF48;    16'd8163: out <= 16'hFDC1;
    16'd8164: out <= 16'hF858;    16'd8165: out <= 16'h02A9;    16'd8166: out <= 16'h01B6;    16'd8167: out <= 16'hFEF0;
    16'd8168: out <= 16'h01AE;    16'd8169: out <= 16'h02C0;    16'd8170: out <= 16'hFDC1;    16'd8171: out <= 16'hFFEA;
    16'd8172: out <= 16'hFFF1;    16'd8173: out <= 16'h0724;    16'd8174: out <= 16'h053D;    16'd8175: out <= 16'hFF2B;
    16'd8176: out <= 16'hFDC8;    16'd8177: out <= 16'h021B;    16'd8178: out <= 16'hFC3D;    16'd8179: out <= 16'hFC49;
    16'd8180: out <= 16'hF8ED;    16'd8181: out <= 16'h05C8;    16'd8182: out <= 16'hFEC5;    16'd8183: out <= 16'h0640;
    16'd8184: out <= 16'h041B;    16'd8185: out <= 16'hFF58;    16'd8186: out <= 16'hFF86;    16'd8187: out <= 16'hFBE3;
    16'd8188: out <= 16'hFF0E;    16'd8189: out <= 16'hFC03;    16'd8190: out <= 16'hFF9D;    16'd8191: out <= 16'hFE50;
    16'd8192: out <= 16'hFFA4;    16'd8193: out <= 16'h06A5;    16'd8194: out <= 16'hFE89;    16'd8195: out <= 16'hFE7C;
    16'd8196: out <= 16'h03E5;    16'd8197: out <= 16'h03A9;    16'd8198: out <= 16'hFD8A;    16'd8199: out <= 16'h04DD;
    16'd8200: out <= 16'h0583;    16'd8201: out <= 16'hFF6A;    16'd8202: out <= 16'h04A7;    16'd8203: out <= 16'h014D;
    16'd8204: out <= 16'hFC20;    16'd8205: out <= 16'hFBE5;    16'd8206: out <= 16'h0441;    16'd8207: out <= 16'h01EA;
    16'd8208: out <= 16'h0319;    16'd8209: out <= 16'h066F;    16'd8210: out <= 16'hFF6D;    16'd8211: out <= 16'hFF3D;
    16'd8212: out <= 16'h04D2;    16'd8213: out <= 16'hFF80;    16'd8214: out <= 16'hFCE9;    16'd8215: out <= 16'hFA78;
    16'd8216: out <= 16'h045B;    16'd8217: out <= 16'h0087;    16'd8218: out <= 16'hFF4A;    16'd8219: out <= 16'h038D;
    16'd8220: out <= 16'hFB9A;    16'd8221: out <= 16'h0398;    16'd8222: out <= 16'h0174;    16'd8223: out <= 16'hF8CA;
    16'd8224: out <= 16'hF950;    16'd8225: out <= 16'h020A;    16'd8226: out <= 16'h0889;    16'd8227: out <= 16'h00AB;
    16'd8228: out <= 16'h016E;    16'd8229: out <= 16'hFB47;    16'd8230: out <= 16'hFDB3;    16'd8231: out <= 16'h01E9;
    16'd8232: out <= 16'h0229;    16'd8233: out <= 16'hF937;    16'd8234: out <= 16'h0045;    16'd8235: out <= 16'h0362;
    16'd8236: out <= 16'h043C;    16'd8237: out <= 16'h04A9;    16'd8238: out <= 16'hFDEE;    16'd8239: out <= 16'hFBEE;
    16'd8240: out <= 16'h08DB;    16'd8241: out <= 16'h06A0;    16'd8242: out <= 16'hFFD9;    16'd8243: out <= 16'h0606;
    16'd8244: out <= 16'h07C4;    16'd8245: out <= 16'h0092;    16'd8246: out <= 16'h067F;    16'd8247: out <= 16'h05DA;
    16'd8248: out <= 16'hFE8C;    16'd8249: out <= 16'h0288;    16'd8250: out <= 16'h02B5;    16'd8251: out <= 16'h0687;
    16'd8252: out <= 16'h0B95;    16'd8253: out <= 16'h059A;    16'd8254: out <= 16'h0849;    16'd8255: out <= 16'h02A1;
    16'd8256: out <= 16'h00EE;    16'd8257: out <= 16'h0912;    16'd8258: out <= 16'hFFF4;    16'd8259: out <= 16'hFF12;
    16'd8260: out <= 16'h02F4;    16'd8261: out <= 16'h08B7;    16'd8262: out <= 16'h0243;    16'd8263: out <= 16'h0487;
    16'd8264: out <= 16'h000F;    16'd8265: out <= 16'h0101;    16'd8266: out <= 16'h0D68;    16'd8267: out <= 16'h02DC;
    16'd8268: out <= 16'h01AC;    16'd8269: out <= 16'h066A;    16'd8270: out <= 16'h0156;    16'd8271: out <= 16'h062E;
    16'd8272: out <= 16'hFAB1;    16'd8273: out <= 16'h12DE;    16'd8274: out <= 16'h05E7;    16'd8275: out <= 16'h059D;
    16'd8276: out <= 16'h08BE;    16'd8277: out <= 16'h0001;    16'd8278: out <= 16'h0062;    16'd8279: out <= 16'h05B1;
    16'd8280: out <= 16'h08A1;    16'd8281: out <= 16'h04B4;    16'd8282: out <= 16'h07D1;    16'd8283: out <= 16'h06A5;
    16'd8284: out <= 16'h0B34;    16'd8285: out <= 16'h0168;    16'd8286: out <= 16'h0421;    16'd8287: out <= 16'h03A7;
    16'd8288: out <= 16'h07BF;    16'd8289: out <= 16'h0014;    16'd8290: out <= 16'hFFA0;    16'd8291: out <= 16'h03F0;
    16'd8292: out <= 16'h0294;    16'd8293: out <= 16'h0660;    16'd8294: out <= 16'h07DB;    16'd8295: out <= 16'h07E2;
    16'd8296: out <= 16'hFEFF;    16'd8297: out <= 16'h03A2;    16'd8298: out <= 16'h0244;    16'd8299: out <= 16'h012C;
    16'd8300: out <= 16'h0218;    16'd8301: out <= 16'hFFAD;    16'd8302: out <= 16'h042B;    16'd8303: out <= 16'h088D;
    16'd8304: out <= 16'hFFA7;    16'd8305: out <= 16'h0349;    16'd8306: out <= 16'h0146;    16'd8307: out <= 16'h00C7;
    16'd8308: out <= 16'h0001;    16'd8309: out <= 16'h00D1;    16'd8310: out <= 16'hFF70;    16'd8311: out <= 16'hFFA2;
    16'd8312: out <= 16'h0290;    16'd8313: out <= 16'hFE39;    16'd8314: out <= 16'h07F1;    16'd8315: out <= 16'h033C;
    16'd8316: out <= 16'h0454;    16'd8317: out <= 16'h0A76;    16'd8318: out <= 16'hFA8A;    16'd8319: out <= 16'h07F4;
    16'd8320: out <= 16'h03B8;    16'd8321: out <= 16'hFFA1;    16'd8322: out <= 16'h01A3;    16'd8323: out <= 16'h0865;
    16'd8324: out <= 16'h0A23;    16'd8325: out <= 16'h0275;    16'd8326: out <= 16'h091E;    16'd8327: out <= 16'hFC0F;
    16'd8328: out <= 16'h051E;    16'd8329: out <= 16'h096F;    16'd8330: out <= 16'h03DE;    16'd8331: out <= 16'h006C;
    16'd8332: out <= 16'h01E5;    16'd8333: out <= 16'h04C7;    16'd8334: out <= 16'h031C;    16'd8335: out <= 16'h041C;
    16'd8336: out <= 16'h0857;    16'd8337: out <= 16'h01B3;    16'd8338: out <= 16'h0221;    16'd8339: out <= 16'h04BF;
    16'd8340: out <= 16'h088E;    16'd8341: out <= 16'h04A7;    16'd8342: out <= 16'h01AA;    16'd8343: out <= 16'hFFA5;
    16'd8344: out <= 16'hFEBD;    16'd8345: out <= 16'h038A;    16'd8346: out <= 16'h037B;    16'd8347: out <= 16'h0781;
    16'd8348: out <= 16'h0A9F;    16'd8349: out <= 16'h05F6;    16'd8350: out <= 16'h0A10;    16'd8351: out <= 16'h0552;
    16'd8352: out <= 16'h0575;    16'd8353: out <= 16'h067A;    16'd8354: out <= 16'hFBE8;    16'd8355: out <= 16'h0659;
    16'd8356: out <= 16'h00EE;    16'd8357: out <= 16'h007E;    16'd8358: out <= 16'h0CB2;    16'd8359: out <= 16'h02F9;
    16'd8360: out <= 16'h0224;    16'd8361: out <= 16'h023A;    16'd8362: out <= 16'h0DF0;    16'd8363: out <= 16'h0A3C;
    16'd8364: out <= 16'h0EFB;    16'd8365: out <= 16'h0636;    16'd8366: out <= 16'h071E;    16'd8367: out <= 16'h0587;
    16'd8368: out <= 16'h0371;    16'd8369: out <= 16'h0506;    16'd8370: out <= 16'h067B;    16'd8371: out <= 16'h01B1;
    16'd8372: out <= 16'h03B8;    16'd8373: out <= 16'h004A;    16'd8374: out <= 16'h0239;    16'd8375: out <= 16'h05EF;
    16'd8376: out <= 16'h09F5;    16'd8377: out <= 16'h06A2;    16'd8378: out <= 16'h0632;    16'd8379: out <= 16'h0952;
    16'd8380: out <= 16'h05FC;    16'd8381: out <= 16'h0220;    16'd8382: out <= 16'h030D;    16'd8383: out <= 16'hFFB2;
    16'd8384: out <= 16'h04CA;    16'd8385: out <= 16'h04A1;    16'd8386: out <= 16'h0BCF;    16'd8387: out <= 16'hFFE8;
    16'd8388: out <= 16'h01C4;    16'd8389: out <= 16'h0502;    16'd8390: out <= 16'h0343;    16'd8391: out <= 16'h0463;
    16'd8392: out <= 16'h0CE8;    16'd8393: out <= 16'h05CB;    16'd8394: out <= 16'h03EC;    16'd8395: out <= 16'hFDC4;
    16'd8396: out <= 16'h00B5;    16'd8397: out <= 16'h01B2;    16'd8398: out <= 16'hFFA7;    16'd8399: out <= 16'h034A;
    16'd8400: out <= 16'hFF55;    16'd8401: out <= 16'h02CC;    16'd8402: out <= 16'h01B3;    16'd8403: out <= 16'hFC56;
    16'd8404: out <= 16'h011C;    16'd8405: out <= 16'hFF58;    16'd8406: out <= 16'h03D0;    16'd8407: out <= 16'hFE19;
    16'd8408: out <= 16'h0035;    16'd8409: out <= 16'h00B8;    16'd8410: out <= 16'hFE58;    16'd8411: out <= 16'hFEAA;
    16'd8412: out <= 16'hFFED;    16'd8413: out <= 16'h00D2;    16'd8414: out <= 16'hFF1F;    16'd8415: out <= 16'hFC58;
    16'd8416: out <= 16'hFD23;    16'd8417: out <= 16'h03DA;    16'd8418: out <= 16'hFC75;    16'd8419: out <= 16'h0492;
    16'd8420: out <= 16'h056A;    16'd8421: out <= 16'hFBB5;    16'd8422: out <= 16'h01CE;    16'd8423: out <= 16'h00F7;
    16'd8424: out <= 16'hFD4A;    16'd8425: out <= 16'hF951;    16'd8426: out <= 16'h04CD;    16'd8427: out <= 16'h0119;
    16'd8428: out <= 16'hFC0E;    16'd8429: out <= 16'hFD39;    16'd8430: out <= 16'hFA43;    16'd8431: out <= 16'hFBDD;
    16'd8432: out <= 16'hFD1E;    16'd8433: out <= 16'h026E;    16'd8434: out <= 16'h0522;    16'd8435: out <= 16'h0061;
    16'd8436: out <= 16'h002B;    16'd8437: out <= 16'h0466;    16'd8438: out <= 16'hFE11;    16'd8439: out <= 16'hFE85;
    16'd8440: out <= 16'h0219;    16'd8441: out <= 16'hFBAF;    16'd8442: out <= 16'hFE4B;    16'd8443: out <= 16'h0000;
    16'd8444: out <= 16'hFC88;    16'd8445: out <= 16'hFE25;    16'd8446: out <= 16'h018B;    16'd8447: out <= 16'hFFC5;
    16'd8448: out <= 16'hFD2F;    16'd8449: out <= 16'h01B0;    16'd8450: out <= 16'hFB5B;    16'd8451: out <= 16'h06E5;
    16'd8452: out <= 16'hFB20;    16'd8453: out <= 16'hFB2D;    16'd8454: out <= 16'h02F0;    16'd8455: out <= 16'h056A;
    16'd8456: out <= 16'hFC1D;    16'd8457: out <= 16'h040E;    16'd8458: out <= 16'hFD66;    16'd8459: out <= 16'h0221;
    16'd8460: out <= 16'h06C2;    16'd8461: out <= 16'hFDA1;    16'd8462: out <= 16'h0131;    16'd8463: out <= 16'h022B;
    16'd8464: out <= 16'h0224;    16'd8465: out <= 16'hFFBF;    16'd8466: out <= 16'hFD61;    16'd8467: out <= 16'hF903;
    16'd8468: out <= 16'hFB25;    16'd8469: out <= 16'h0587;    16'd8470: out <= 16'hFF56;    16'd8471: out <= 16'hFA96;
    16'd8472: out <= 16'hFF70;    16'd8473: out <= 16'h0258;    16'd8474: out <= 16'h03D8;    16'd8475: out <= 16'hFDA7;
    16'd8476: out <= 16'hFBED;    16'd8477: out <= 16'hFD35;    16'd8478: out <= 16'h012C;    16'd8479: out <= 16'hFDBD;
    16'd8480: out <= 16'hFFE7;    16'd8481: out <= 16'h053A;    16'd8482: out <= 16'h04A7;    16'd8483: out <= 16'h00CB;
    16'd8484: out <= 16'h032A;    16'd8485: out <= 16'hFAC5;    16'd8486: out <= 16'hFF8F;    16'd8487: out <= 16'hFBAE;
    16'd8488: out <= 16'hFD94;    16'd8489: out <= 16'h002D;    16'd8490: out <= 16'h0136;    16'd8491: out <= 16'h0297;
    16'd8492: out <= 16'h0552;    16'd8493: out <= 16'h0A30;    16'd8494: out <= 16'h0185;    16'd8495: out <= 16'hFE41;
    16'd8496: out <= 16'h05B7;    16'd8497: out <= 16'h034E;    16'd8498: out <= 16'h0849;    16'd8499: out <= 16'h092B;
    16'd8500: out <= 16'h009E;    16'd8501: out <= 16'h010E;    16'd8502: out <= 16'h0B8C;    16'd8503: out <= 16'h04EA;
    16'd8504: out <= 16'h02EC;    16'd8505: out <= 16'h0497;    16'd8506: out <= 16'h016F;    16'd8507: out <= 16'h00DC;
    16'd8508: out <= 16'h01E1;    16'd8509: out <= 16'h07E6;    16'd8510: out <= 16'h0481;    16'd8511: out <= 16'h0604;
    16'd8512: out <= 16'h0533;    16'd8513: out <= 16'h057F;    16'd8514: out <= 16'h0A37;    16'd8515: out <= 16'h0340;
    16'd8516: out <= 16'h0256;    16'd8517: out <= 16'h0533;    16'd8518: out <= 16'h022C;    16'd8519: out <= 16'h027C;
    16'd8520: out <= 16'h02D2;    16'd8521: out <= 16'hFF65;    16'd8522: out <= 16'hFBA5;    16'd8523: out <= 16'h0038;
    16'd8524: out <= 16'h023C;    16'd8525: out <= 16'h00F6;    16'd8526: out <= 16'hFE70;    16'd8527: out <= 16'h0044;
    16'd8528: out <= 16'h00B4;    16'd8529: out <= 16'hFDFD;    16'd8530: out <= 16'h0339;    16'd8531: out <= 16'h0544;
    16'd8532: out <= 16'hFF43;    16'd8533: out <= 16'hFE78;    16'd8534: out <= 16'h025B;    16'd8535: out <= 16'hFD1F;
    16'd8536: out <= 16'h0372;    16'd8537: out <= 16'hFCC1;    16'd8538: out <= 16'h0882;    16'd8539: out <= 16'h0079;
    16'd8540: out <= 16'h07F6;    16'd8541: out <= 16'h01A9;    16'd8542: out <= 16'h0245;    16'd8543: out <= 16'h039A;
    16'd8544: out <= 16'h01DE;    16'd8545: out <= 16'h080A;    16'd8546: out <= 16'h0467;    16'd8547: out <= 16'h033B;
    16'd8548: out <= 16'h0884;    16'd8549: out <= 16'h08B2;    16'd8550: out <= 16'h00BC;    16'd8551: out <= 16'h0507;
    16'd8552: out <= 16'h0662;    16'd8553: out <= 16'h05EF;    16'd8554: out <= 16'h01B1;    16'd8555: out <= 16'hFF83;
    16'd8556: out <= 16'hFE1A;    16'd8557: out <= 16'h04B2;    16'd8558: out <= 16'h05D9;    16'd8559: out <= 16'hFE74;
    16'd8560: out <= 16'h0726;    16'd8561: out <= 16'h0B60;    16'd8562: out <= 16'h0498;    16'd8563: out <= 16'h0A00;
    16'd8564: out <= 16'h0206;    16'd8565: out <= 16'h0837;    16'd8566: out <= 16'h058C;    16'd8567: out <= 16'hFEB1;
    16'd8568: out <= 16'h02B3;    16'd8569: out <= 16'h05A7;    16'd8570: out <= 16'h06DD;    16'd8571: out <= 16'h052C;
    16'd8572: out <= 16'h082B;    16'd8573: out <= 16'h0296;    16'd8574: out <= 16'hFC2A;    16'd8575: out <= 16'h02F0;
    16'd8576: out <= 16'h01B3;    16'd8577: out <= 16'h0828;    16'd8578: out <= 16'h03F6;    16'd8579: out <= 16'hFF76;
    16'd8580: out <= 16'h08BB;    16'd8581: out <= 16'h02A0;    16'd8582: out <= 16'h0BEE;    16'd8583: out <= 16'h086F;
    16'd8584: out <= 16'hFFCC;    16'd8585: out <= 16'h0575;    16'd8586: out <= 16'h030B;    16'd8587: out <= 16'h064B;
    16'd8588: out <= 16'hFB12;    16'd8589: out <= 16'h07A3;    16'd8590: out <= 16'hFEDB;    16'd8591: out <= 16'hFE70;
    16'd8592: out <= 16'h0450;    16'd8593: out <= 16'h0617;    16'd8594: out <= 16'h0258;    16'd8595: out <= 16'h07C0;
    16'd8596: out <= 16'h060F;    16'd8597: out <= 16'h086C;    16'd8598: out <= 16'h0877;    16'd8599: out <= 16'h0477;
    16'd8600: out <= 16'h0406;    16'd8601: out <= 16'h02A8;    16'd8602: out <= 16'h03B3;    16'd8603: out <= 16'hFFAA;
    16'd8604: out <= 16'h022F;    16'd8605: out <= 16'h058E;    16'd8606: out <= 16'h0567;    16'd8607: out <= 16'h01DB;
    16'd8608: out <= 16'h05E7;    16'd8609: out <= 16'h0024;    16'd8610: out <= 16'h0100;    16'd8611: out <= 16'h053A;
    16'd8612: out <= 16'hFC78;    16'd8613: out <= 16'h0A9D;    16'd8614: out <= 16'h05D5;    16'd8615: out <= 16'hFC45;
    16'd8616: out <= 16'h0AD5;    16'd8617: out <= 16'hFD6B;    16'd8618: out <= 16'h0773;    16'd8619: out <= 16'h091C;
    16'd8620: out <= 16'h03E7;    16'd8621: out <= 16'h0390;    16'd8622: out <= 16'hF874;    16'd8623: out <= 16'h0464;
    16'd8624: out <= 16'hFB7F;    16'd8625: out <= 16'h003E;    16'd8626: out <= 16'h082B;    16'd8627: out <= 16'h0714;
    16'd8628: out <= 16'hFDC2;    16'd8629: out <= 16'h0126;    16'd8630: out <= 16'h0786;    16'd8631: out <= 16'hFEA4;
    16'd8632: out <= 16'h03D6;    16'd8633: out <= 16'h0125;    16'd8634: out <= 16'h0ADA;    16'd8635: out <= 16'h0310;
    16'd8636: out <= 16'h0B5E;    16'd8637: out <= 16'h0783;    16'd8638: out <= 16'h00F0;    16'd8639: out <= 16'h04F6;
    16'd8640: out <= 16'h0600;    16'd8641: out <= 16'hFC0A;    16'd8642: out <= 16'h0A7D;    16'd8643: out <= 16'h0185;
    16'd8644: out <= 16'h002A;    16'd8645: out <= 16'hFDA1;    16'd8646: out <= 16'hF9BF;    16'd8647: out <= 16'h00E9;
    16'd8648: out <= 16'h02C2;    16'd8649: out <= 16'h0497;    16'd8650: out <= 16'h0CD4;    16'd8651: out <= 16'hFF5E;
    16'd8652: out <= 16'h02C3;    16'd8653: out <= 16'hFEC7;    16'd8654: out <= 16'hFF30;    16'd8655: out <= 16'hF86F;
    16'd8656: out <= 16'hFEAD;    16'd8657: out <= 16'hFF19;    16'd8658: out <= 16'hFED3;    16'd8659: out <= 16'hFFAE;
    16'd8660: out <= 16'hFA74;    16'd8661: out <= 16'h00C9;    16'd8662: out <= 16'hFCDD;    16'd8663: out <= 16'hFF05;
    16'd8664: out <= 16'hFDC6;    16'd8665: out <= 16'h0604;    16'd8666: out <= 16'hFF21;    16'd8667: out <= 16'hF7CA;
    16'd8668: out <= 16'hFAEA;    16'd8669: out <= 16'h02F1;    16'd8670: out <= 16'hFFB3;    16'd8671: out <= 16'hFD20;
    16'd8672: out <= 16'hFD4B;    16'd8673: out <= 16'hFA47;    16'd8674: out <= 16'h01F6;    16'd8675: out <= 16'hFE41;
    16'd8676: out <= 16'h038F;    16'd8677: out <= 16'hFEC6;    16'd8678: out <= 16'h024B;    16'd8679: out <= 16'hFF5B;
    16'd8680: out <= 16'h02B5;    16'd8681: out <= 16'h014B;    16'd8682: out <= 16'hFE60;    16'd8683: out <= 16'hFEA4;
    16'd8684: out <= 16'h0401;    16'd8685: out <= 16'h0013;    16'd8686: out <= 16'hFD52;    16'd8687: out <= 16'hFDA8;
    16'd8688: out <= 16'hFDBF;    16'd8689: out <= 16'hFFBF;    16'd8690: out <= 16'hFFAE;    16'd8691: out <= 16'hFFB6;
    16'd8692: out <= 16'hFCA2;    16'd8693: out <= 16'hFB7A;    16'd8694: out <= 16'h08E4;    16'd8695: out <= 16'h0054;
    16'd8696: out <= 16'h031B;    16'd8697: out <= 16'hFD30;    16'd8698: out <= 16'hFF76;    16'd8699: out <= 16'hFD62;
    16'd8700: out <= 16'h0142;    16'd8701: out <= 16'hFDEF;    16'd8702: out <= 16'hF9E4;    16'd8703: out <= 16'h00EA;
    16'd8704: out <= 16'h03C7;    16'd8705: out <= 16'hFD61;    16'd8706: out <= 16'h0091;    16'd8707: out <= 16'hF728;
    16'd8708: out <= 16'h0313;    16'd8709: out <= 16'h00C2;    16'd8710: out <= 16'h0094;    16'd8711: out <= 16'hFEF5;
    16'd8712: out <= 16'hFE65;    16'd8713: out <= 16'hFE43;    16'd8714: out <= 16'hF9EB;    16'd8715: out <= 16'h01FD;
    16'd8716: out <= 16'h0439;    16'd8717: out <= 16'hFECE;    16'd8718: out <= 16'h00F4;    16'd8719: out <= 16'hFCE6;
    16'd8720: out <= 16'hFB24;    16'd8721: out <= 16'hFD1D;    16'd8722: out <= 16'h037F;    16'd8723: out <= 16'hFE88;
    16'd8724: out <= 16'h0176;    16'd8725: out <= 16'hFD29;    16'd8726: out <= 16'h0240;    16'd8727: out <= 16'h008D;
    16'd8728: out <= 16'hFFBB;    16'd8729: out <= 16'hFE7C;    16'd8730: out <= 16'h05BC;    16'd8731: out <= 16'h01E9;
    16'd8732: out <= 16'h0101;    16'd8733: out <= 16'h02E7;    16'd8734: out <= 16'h00A9;    16'd8735: out <= 16'h034E;
    16'd8736: out <= 16'hFF4E;    16'd8737: out <= 16'h006A;    16'd8738: out <= 16'h06D5;    16'd8739: out <= 16'h01F8;
    16'd8740: out <= 16'h0613;    16'd8741: out <= 16'h0473;    16'd8742: out <= 16'hF8F1;    16'd8743: out <= 16'h04E3;
    16'd8744: out <= 16'h04E3;    16'd8745: out <= 16'h0110;    16'd8746: out <= 16'h05B6;    16'd8747: out <= 16'hFD17;
    16'd8748: out <= 16'h06C1;    16'd8749: out <= 16'hFA65;    16'd8750: out <= 16'hFCCC;    16'd8751: out <= 16'h00A4;
    16'd8752: out <= 16'h044F;    16'd8753: out <= 16'h0148;    16'd8754: out <= 16'h05A6;    16'd8755: out <= 16'h04FB;
    16'd8756: out <= 16'h052A;    16'd8757: out <= 16'h07BE;    16'd8758: out <= 16'h05EE;    16'd8759: out <= 16'h0989;
    16'd8760: out <= 16'h01C8;    16'd8761: out <= 16'h08A4;    16'd8762: out <= 16'h067C;    16'd8763: out <= 16'h0233;
    16'd8764: out <= 16'h04D1;    16'd8765: out <= 16'h093F;    16'd8766: out <= 16'h051E;    16'd8767: out <= 16'h0223;
    16'd8768: out <= 16'h057B;    16'd8769: out <= 16'hFE13;    16'd8770: out <= 16'h038A;    16'd8771: out <= 16'h01CC;
    16'd8772: out <= 16'h0322;    16'd8773: out <= 16'h082B;    16'd8774: out <= 16'h010A;    16'd8775: out <= 16'hFFD8;
    16'd8776: out <= 16'h0210;    16'd8777: out <= 16'h02E6;    16'd8778: out <= 16'h029E;    16'd8779: out <= 16'h0125;
    16'd8780: out <= 16'h0BD5;    16'd8781: out <= 16'h06DA;    16'd8782: out <= 16'h05EA;    16'd8783: out <= 16'h044D;
    16'd8784: out <= 16'h01FA;    16'd8785: out <= 16'h0730;    16'd8786: out <= 16'h10A8;    16'd8787: out <= 16'h060F;
    16'd8788: out <= 16'h02A6;    16'd8789: out <= 16'h0359;    16'd8790: out <= 16'h08D1;    16'd8791: out <= 16'h00FD;
    16'd8792: out <= 16'h065E;    16'd8793: out <= 16'h0457;    16'd8794: out <= 16'h0442;    16'd8795: out <= 16'h01DD;
    16'd8796: out <= 16'h05A9;    16'd8797: out <= 16'h0624;    16'd8798: out <= 16'h0254;    16'd8799: out <= 16'h0710;
    16'd8800: out <= 16'h03E1;    16'd8801: out <= 16'h059D;    16'd8802: out <= 16'hFD9F;    16'd8803: out <= 16'h0611;
    16'd8804: out <= 16'h03BC;    16'd8805: out <= 16'h03DA;    16'd8806: out <= 16'h05A8;    16'd8807: out <= 16'hFEF6;
    16'd8808: out <= 16'h0B36;    16'd8809: out <= 16'h0081;    16'd8810: out <= 16'h0913;    16'd8811: out <= 16'h02A3;
    16'd8812: out <= 16'h0D48;    16'd8813: out <= 16'h0986;    16'd8814: out <= 16'h00FC;    16'd8815: out <= 16'h037F;
    16'd8816: out <= 16'h0422;    16'd8817: out <= 16'h05EF;    16'd8818: out <= 16'hFE54;    16'd8819: out <= 16'h00AE;
    16'd8820: out <= 16'h042A;    16'd8821: out <= 16'h03DC;    16'd8822: out <= 16'h0843;    16'd8823: out <= 16'h02EB;
    16'd8824: out <= 16'h02E7;    16'd8825: out <= 16'h083F;    16'd8826: out <= 16'hFFF8;    16'd8827: out <= 16'hFBFE;
    16'd8828: out <= 16'h01A4;    16'd8829: out <= 16'h024C;    16'd8830: out <= 16'h05DC;    16'd8831: out <= 16'h0694;
    16'd8832: out <= 16'h0485;    16'd8833: out <= 16'h050B;    16'd8834: out <= 16'hFA3C;    16'd8835: out <= 16'hFD95;
    16'd8836: out <= 16'h0711;    16'd8837: out <= 16'h058D;    16'd8838: out <= 16'h0742;    16'd8839: out <= 16'hFF8E;
    16'd8840: out <= 16'h093F;    16'd8841: out <= 16'h070B;    16'd8842: out <= 16'h059D;    16'd8843: out <= 16'hFE95;
    16'd8844: out <= 16'h03C7;    16'd8845: out <= 16'hFC7A;    16'd8846: out <= 16'hFA23;    16'd8847: out <= 16'hFE58;
    16'd8848: out <= 16'h0898;    16'd8849: out <= 16'h00A4;    16'd8850: out <= 16'h0450;    16'd8851: out <= 16'h03EB;
    16'd8852: out <= 16'h05EA;    16'd8853: out <= 16'h038E;    16'd8854: out <= 16'h06DD;    16'd8855: out <= 16'h03E6;
    16'd8856: out <= 16'h02A5;    16'd8857: out <= 16'h00E8;    16'd8858: out <= 16'hFE7F;    16'd8859: out <= 16'h083E;
    16'd8860: out <= 16'hFFA3;    16'd8861: out <= 16'h02EF;    16'd8862: out <= 16'h0547;    16'd8863: out <= 16'h0268;
    16'd8864: out <= 16'hFA0B;    16'd8865: out <= 16'h05F6;    16'd8866: out <= 16'h05A6;    16'd8867: out <= 16'hFF7B;
    16'd8868: out <= 16'h081A;    16'd8869: out <= 16'hFF28;    16'd8870: out <= 16'h04B5;    16'd8871: out <= 16'h09C4;
    16'd8872: out <= 16'h0527;    16'd8873: out <= 16'h0673;    16'd8874: out <= 16'h093C;    16'd8875: out <= 16'h06C1;
    16'd8876: out <= 16'h02A4;    16'd8877: out <= 16'h02BF;    16'd8878: out <= 16'hFE49;    16'd8879: out <= 16'hFBF3;
    16'd8880: out <= 16'h04FE;    16'd8881: out <= 16'hFEE7;    16'd8882: out <= 16'h0884;    16'd8883: out <= 16'h07C2;
    16'd8884: out <= 16'h09B2;    16'd8885: out <= 16'h02A2;    16'd8886: out <= 16'h0538;    16'd8887: out <= 16'h09C3;
    16'd8888: out <= 16'h0A9B;    16'd8889: out <= 16'h02A3;    16'd8890: out <= 16'h0258;    16'd8891: out <= 16'hFEFD;
    16'd8892: out <= 16'h0760;    16'd8893: out <= 16'h0115;    16'd8894: out <= 16'h05B8;    16'd8895: out <= 16'h066B;
    16'd8896: out <= 16'h0487;    16'd8897: out <= 16'h0CD9;    16'd8898: out <= 16'h04DB;    16'd8899: out <= 16'h05C9;
    16'd8900: out <= 16'h049F;    16'd8901: out <= 16'h0A48;    16'd8902: out <= 16'h04FD;    16'd8903: out <= 16'h0013;
    16'd8904: out <= 16'h0804;    16'd8905: out <= 16'h05DB;    16'd8906: out <= 16'h007B;    16'd8907: out <= 16'h055D;
    16'd8908: out <= 16'hFF57;    16'd8909: out <= 16'h0451;    16'd8910: out <= 16'hFD3C;    16'd8911: out <= 16'h00B7;
    16'd8912: out <= 16'hF985;    16'd8913: out <= 16'hFD02;    16'd8914: out <= 16'h0239;    16'd8915: out <= 16'h054C;
    16'd8916: out <= 16'h0497;    16'd8917: out <= 16'hFFF1;    16'd8918: out <= 16'hFFA1;    16'd8919: out <= 16'h01B1;
    16'd8920: out <= 16'h05BE;    16'd8921: out <= 16'hFFEB;    16'd8922: out <= 16'hFC95;    16'd8923: out <= 16'hFDA5;
    16'd8924: out <= 16'hFD22;    16'd8925: out <= 16'hFF03;    16'd8926: out <= 16'h02A1;    16'd8927: out <= 16'h04F6;
    16'd8928: out <= 16'hFFB8;    16'd8929: out <= 16'hFEA2;    16'd8930: out <= 16'hF97E;    16'd8931: out <= 16'h026E;
    16'd8932: out <= 16'h003A;    16'd8933: out <= 16'hFE56;    16'd8934: out <= 16'hF7DA;    16'd8935: out <= 16'hFB43;
    16'd8936: out <= 16'hFCE5;    16'd8937: out <= 16'h00D7;    16'd8938: out <= 16'hFF25;    16'd8939: out <= 16'h094E;
    16'd8940: out <= 16'hFF80;    16'd8941: out <= 16'h021D;    16'd8942: out <= 16'h0816;    16'd8943: out <= 16'hFE90;
    16'd8944: out <= 16'hF7B8;    16'd8945: out <= 16'hFE42;    16'd8946: out <= 16'h0621;    16'd8947: out <= 16'hFDB7;
    16'd8948: out <= 16'h05B8;    16'd8949: out <= 16'h007F;    16'd8950: out <= 16'h0398;    16'd8951: out <= 16'h0734;
    16'd8952: out <= 16'h02BB;    16'd8953: out <= 16'h01C9;    16'd8954: out <= 16'hFF72;    16'd8955: out <= 16'hFF91;
    16'd8956: out <= 16'h0083;    16'd8957: out <= 16'hFEE4;    16'd8958: out <= 16'hFFFA;    16'd8959: out <= 16'hFA31;
    16'd8960: out <= 16'hFB87;    16'd8961: out <= 16'hFD36;    16'd8962: out <= 16'h0A8F;    16'd8963: out <= 16'h02C5;
    16'd8964: out <= 16'h04FA;    16'd8965: out <= 16'hFEC6;    16'd8966: out <= 16'hFE00;    16'd8967: out <= 16'hFCAE;
    16'd8968: out <= 16'hFD40;    16'd8969: out <= 16'hFDB2;    16'd8970: out <= 16'hF92A;    16'd8971: out <= 16'h02FA;
    16'd8972: out <= 16'h0573;    16'd8973: out <= 16'h02F7;    16'd8974: out <= 16'hF8EC;    16'd8975: out <= 16'h0204;
    16'd8976: out <= 16'h013B;    16'd8977: out <= 16'h018E;    16'd8978: out <= 16'hFD11;    16'd8979: out <= 16'h074E;
    16'd8980: out <= 16'h024F;    16'd8981: out <= 16'hF593;    16'd8982: out <= 16'hFEAC;    16'd8983: out <= 16'hFCC2;
    16'd8984: out <= 16'hFA3B;    16'd8985: out <= 16'hFA09;    16'd8986: out <= 16'hFCB0;    16'd8987: out <= 16'hF9F1;
    16'd8988: out <= 16'h023E;    16'd8989: out <= 16'hFD09;    16'd8990: out <= 16'hFFF8;    16'd8991: out <= 16'h055B;
    16'd8992: out <= 16'h0347;    16'd8993: out <= 16'hFFAA;    16'd8994: out <= 16'h0117;    16'd8995: out <= 16'h0337;
    16'd8996: out <= 16'hFD83;    16'd8997: out <= 16'h003D;    16'd8998: out <= 16'h059F;    16'd8999: out <= 16'h0338;
    16'd9000: out <= 16'h0867;    16'd9001: out <= 16'h08EC;    16'd9002: out <= 16'hFF1A;    16'd9003: out <= 16'hFC3B;
    16'd9004: out <= 16'hF81B;    16'd9005: out <= 16'hFE94;    16'd9006: out <= 16'h01FA;    16'd9007: out <= 16'h0266;
    16'd9008: out <= 16'h044F;    16'd9009: out <= 16'h0264;    16'd9010: out <= 16'h051D;    16'd9011: out <= 16'h0470;
    16'd9012: out <= 16'h089A;    16'd9013: out <= 16'h04EB;    16'd9014: out <= 16'h0494;    16'd9015: out <= 16'h04E2;
    16'd9016: out <= 16'h0085;    16'd9017: out <= 16'h0861;    16'd9018: out <= 16'h00CB;    16'd9019: out <= 16'hFFDC;
    16'd9020: out <= 16'h06D6;    16'd9021: out <= 16'h057E;    16'd9022: out <= 16'h01A4;    16'd9023: out <= 16'h002C;
    16'd9024: out <= 16'h0317;    16'd9025: out <= 16'h024B;    16'd9026: out <= 16'h0976;    16'd9027: out <= 16'h06F6;
    16'd9028: out <= 16'h0A50;    16'd9029: out <= 16'hFCB0;    16'd9030: out <= 16'hFED1;    16'd9031: out <= 16'h058C;
    16'd9032: out <= 16'h0D5B;    16'd9033: out <= 16'h0663;    16'd9034: out <= 16'h0282;    16'd9035: out <= 16'h0868;
    16'd9036: out <= 16'h0201;    16'd9037: out <= 16'h0259;    16'd9038: out <= 16'hFB7B;    16'd9039: out <= 16'h0894;
    16'd9040: out <= 16'h03C6;    16'd9041: out <= 16'h07FE;    16'd9042: out <= 16'h0640;    16'd9043: out <= 16'h04E1;
    16'd9044: out <= 16'h0270;    16'd9045: out <= 16'hFDA8;    16'd9046: out <= 16'h04CB;    16'd9047: out <= 16'h02F7;
    16'd9048: out <= 16'h01C0;    16'd9049: out <= 16'h0029;    16'd9050: out <= 16'h08CF;    16'd9051: out <= 16'hFF4C;
    16'd9052: out <= 16'h0798;    16'd9053: out <= 16'hFFCE;    16'd9054: out <= 16'h061C;    16'd9055: out <= 16'h01F7;
    16'd9056: out <= 16'h0556;    16'd9057: out <= 16'h023E;    16'd9058: out <= 16'h0A05;    16'd9059: out <= 16'h0518;
    16'd9060: out <= 16'h0682;    16'd9061: out <= 16'h092C;    16'd9062: out <= 16'hFD26;    16'd9063: out <= 16'h0372;
    16'd9064: out <= 16'h03A8;    16'd9065: out <= 16'hFE5C;    16'd9066: out <= 16'h02A9;    16'd9067: out <= 16'h0470;
    16'd9068: out <= 16'h0364;    16'd9069: out <= 16'h0808;    16'd9070: out <= 16'h067D;    16'd9071: out <= 16'h0210;
    16'd9072: out <= 16'h094E;    16'd9073: out <= 16'h0383;    16'd9074: out <= 16'h016F;    16'd9075: out <= 16'h0126;
    16'd9076: out <= 16'h0409;    16'd9077: out <= 16'hFFB3;    16'd9078: out <= 16'hFF73;    16'd9079: out <= 16'hFC40;
    16'd9080: out <= 16'h029A;    16'd9081: out <= 16'hFE69;    16'd9082: out <= 16'h0110;    16'd9083: out <= 16'h05DF;
    16'd9084: out <= 16'h06CE;    16'd9085: out <= 16'h039D;    16'd9086: out <= 16'h06BE;    16'd9087: out <= 16'hFD16;
    16'd9088: out <= 16'h0BC4;    16'd9089: out <= 16'h066E;    16'd9090: out <= 16'h03C9;    16'd9091: out <= 16'h0497;
    16'd9092: out <= 16'h08B4;    16'd9093: out <= 16'h03BA;    16'd9094: out <= 16'h05FE;    16'd9095: out <= 16'h0605;
    16'd9096: out <= 16'h051D;    16'd9097: out <= 16'h052D;    16'd9098: out <= 16'h07EF;    16'd9099: out <= 16'h0060;
    16'd9100: out <= 16'h08BF;    16'd9101: out <= 16'h0315;    16'd9102: out <= 16'h09D4;    16'd9103: out <= 16'hFFCC;
    16'd9104: out <= 16'h0729;    16'd9105: out <= 16'hFFD0;    16'd9106: out <= 16'hFF9B;    16'd9107: out <= 16'hFED3;
    16'd9108: out <= 16'h0425;    16'd9109: out <= 16'h05B7;    16'd9110: out <= 16'hFECC;    16'd9111: out <= 16'h076B;
    16'd9112: out <= 16'hFEC8;    16'd9113: out <= 16'h0695;    16'd9114: out <= 16'hFF80;    16'd9115: out <= 16'hFD6E;
    16'd9116: out <= 16'h07A0;    16'd9117: out <= 16'h0263;    16'd9118: out <= 16'h0467;    16'd9119: out <= 16'h0569;
    16'd9120: out <= 16'h027C;    16'd9121: out <= 16'hFFE3;    16'd9122: out <= 16'h0019;    16'd9123: out <= 16'h026A;
    16'd9124: out <= 16'h051F;    16'd9125: out <= 16'h0A48;    16'd9126: out <= 16'h071F;    16'd9127: out <= 16'h002B;
    16'd9128: out <= 16'h079F;    16'd9129: out <= 16'hFDC4;    16'd9130: out <= 16'hFDB6;    16'd9131: out <= 16'h053E;
    16'd9132: out <= 16'h01B8;    16'd9133: out <= 16'h01E6;    16'd9134: out <= 16'h0181;    16'd9135: out <= 16'h0672;
    16'd9136: out <= 16'h04FE;    16'd9137: out <= 16'h0A41;    16'd9138: out <= 16'h0643;    16'd9139: out <= 16'hFF04;
    16'd9140: out <= 16'hFF15;    16'd9141: out <= 16'hFC96;    16'd9142: out <= 16'h0378;    16'd9143: out <= 16'h0BEF;
    16'd9144: out <= 16'h02A4;    16'd9145: out <= 16'hFF4B;    16'd9146: out <= 16'h06EF;    16'd9147: out <= 16'h0090;
    16'd9148: out <= 16'hFF82;    16'd9149: out <= 16'h06A2;    16'd9150: out <= 16'h0A16;    16'd9151: out <= 16'hFE91;
    16'd9152: out <= 16'hFD37;    16'd9153: out <= 16'h0202;    16'd9154: out <= 16'h0635;    16'd9155: out <= 16'h0810;
    16'd9156: out <= 16'hFF5D;    16'd9157: out <= 16'h0BEE;    16'd9158: out <= 16'h04D6;    16'd9159: out <= 16'hFF1F;
    16'd9160: out <= 16'h0991;    16'd9161: out <= 16'h036D;    16'd9162: out <= 16'h01DD;    16'd9163: out <= 16'h04BC;
    16'd9164: out <= 16'h0274;    16'd9165: out <= 16'hFCA4;    16'd9166: out <= 16'hF992;    16'd9167: out <= 16'hFCF8;
    16'd9168: out <= 16'h0321;    16'd9169: out <= 16'h0043;    16'd9170: out <= 16'h0086;    16'd9171: out <= 16'h07B2;
    16'd9172: out <= 16'hFB8B;    16'd9173: out <= 16'h0209;    16'd9174: out <= 16'h017C;    16'd9175: out <= 16'hFFF6;
    16'd9176: out <= 16'h0557;    16'd9177: out <= 16'h0616;    16'd9178: out <= 16'h0147;    16'd9179: out <= 16'hFF80;
    16'd9180: out <= 16'h038D;    16'd9181: out <= 16'h0334;    16'd9182: out <= 16'h06A4;    16'd9183: out <= 16'h0B16;
    16'd9184: out <= 16'h086F;    16'd9185: out <= 16'hFCFE;    16'd9186: out <= 16'h01B9;    16'd9187: out <= 16'h03AA;
    16'd9188: out <= 16'hFD0F;    16'd9189: out <= 16'h03D0;    16'd9190: out <= 16'h0283;    16'd9191: out <= 16'h0061;
    16'd9192: out <= 16'h02F0;    16'd9193: out <= 16'hFC85;    16'd9194: out <= 16'h0005;    16'd9195: out <= 16'h0073;
    16'd9196: out <= 16'h0267;    16'd9197: out <= 16'h070D;    16'd9198: out <= 16'h00E5;    16'd9199: out <= 16'hFFD6;
    16'd9200: out <= 16'h0089;    16'd9201: out <= 16'h0039;    16'd9202: out <= 16'h0154;    16'd9203: out <= 16'hF944;
    16'd9204: out <= 16'hFF4D;    16'd9205: out <= 16'hFF51;    16'd9206: out <= 16'hFB68;    16'd9207: out <= 16'h051B;
    16'd9208: out <= 16'hF8DF;    16'd9209: out <= 16'hFB49;    16'd9210: out <= 16'h00D2;    16'd9211: out <= 16'hFDF4;
    16'd9212: out <= 16'hF891;    16'd9213: out <= 16'h0251;    16'd9214: out <= 16'h0491;    16'd9215: out <= 16'hFDC4;
    16'd9216: out <= 16'h0429;    16'd9217: out <= 16'h0568;    16'd9218: out <= 16'hFAA1;    16'd9219: out <= 16'h021B;
    16'd9220: out <= 16'h00C0;    16'd9221: out <= 16'h06B0;    16'd9222: out <= 16'h02B8;    16'd9223: out <= 16'hFED0;
    16'd9224: out <= 16'h0342;    16'd9225: out <= 16'hFCD9;    16'd9226: out <= 16'hFF52;    16'd9227: out <= 16'hFE48;
    16'd9228: out <= 16'h00C9;    16'd9229: out <= 16'hFD75;    16'd9230: out <= 16'h0977;    16'd9231: out <= 16'hFEBD;
    16'd9232: out <= 16'h03B3;    16'd9233: out <= 16'hFD20;    16'd9234: out <= 16'hF875;    16'd9235: out <= 16'hFE2B;
    16'd9236: out <= 16'hFE4D;    16'd9237: out <= 16'h00AD;    16'd9238: out <= 16'h00E4;    16'd9239: out <= 16'h060A;
    16'd9240: out <= 16'hF816;    16'd9241: out <= 16'hFF9E;    16'd9242: out <= 16'h0441;    16'd9243: out <= 16'hF971;
    16'd9244: out <= 16'h02E2;    16'd9245: out <= 16'h01DC;    16'd9246: out <= 16'hFB61;    16'd9247: out <= 16'h0065;
    16'd9248: out <= 16'hFE56;    16'd9249: out <= 16'hFE43;    16'd9250: out <= 16'h0067;    16'd9251: out <= 16'hFC89;
    16'd9252: out <= 16'hF87C;    16'd9253: out <= 16'h0399;    16'd9254: out <= 16'h04D4;    16'd9255: out <= 16'h0825;
    16'd9256: out <= 16'h02EE;    16'd9257: out <= 16'h0678;    16'd9258: out <= 16'hFBF4;    16'd9259: out <= 16'h02F5;
    16'd9260: out <= 16'hFC69;    16'd9261: out <= 16'hFE4E;    16'd9262: out <= 16'h0452;    16'd9263: out <= 16'hFF8A;
    16'd9264: out <= 16'h051F;    16'd9265: out <= 16'hFEA2;    16'd9266: out <= 16'h0286;    16'd9267: out <= 16'h074D;
    16'd9268: out <= 16'h03AD;    16'd9269: out <= 16'h059C;    16'd9270: out <= 16'h035F;    16'd9271: out <= 16'h023F;
    16'd9272: out <= 16'h07D5;    16'd9273: out <= 16'h071B;    16'd9274: out <= 16'hFF69;    16'd9275: out <= 16'h0218;
    16'd9276: out <= 16'h02A6;    16'd9277: out <= 16'h0708;    16'd9278: out <= 16'h04CE;    16'd9279: out <= 16'h0083;
    16'd9280: out <= 16'h0290;    16'd9281: out <= 16'h033E;    16'd9282: out <= 16'h052C;    16'd9283: out <= 16'h04E2;
    16'd9284: out <= 16'hFE7F;    16'd9285: out <= 16'h05B7;    16'd9286: out <= 16'h00F2;    16'd9287: out <= 16'h08A5;
    16'd9288: out <= 16'hFEB6;    16'd9289: out <= 16'h069E;    16'd9290: out <= 16'h0D8C;    16'd9291: out <= 16'h01E0;
    16'd9292: out <= 16'h08D1;    16'd9293: out <= 16'h04C9;    16'd9294: out <= 16'h0B13;    16'd9295: out <= 16'h031F;
    16'd9296: out <= 16'h035B;    16'd9297: out <= 16'h088B;    16'd9298: out <= 16'h0218;    16'd9299: out <= 16'h07FC;
    16'd9300: out <= 16'hFF3A;    16'd9301: out <= 16'h0AC9;    16'd9302: out <= 16'hF9AC;    16'd9303: out <= 16'h022A;
    16'd9304: out <= 16'h0A97;    16'd9305: out <= 16'h0B93;    16'd9306: out <= 16'h027A;    16'd9307: out <= 16'h0575;
    16'd9308: out <= 16'h06DF;    16'd9309: out <= 16'hFFA0;    16'd9310: out <= 16'h0332;    16'd9311: out <= 16'h0871;
    16'd9312: out <= 16'h02B2;    16'd9313: out <= 16'h0651;    16'd9314: out <= 16'h0BF0;    16'd9315: out <= 16'h008D;
    16'd9316: out <= 16'h0896;    16'd9317: out <= 16'h06F8;    16'd9318: out <= 16'h04A1;    16'd9319: out <= 16'h0432;
    16'd9320: out <= 16'h063F;    16'd9321: out <= 16'h0377;    16'd9322: out <= 16'h02F4;    16'd9323: out <= 16'h02C6;
    16'd9324: out <= 16'h0015;    16'd9325: out <= 16'h081D;    16'd9326: out <= 16'h07A5;    16'd9327: out <= 16'h0038;
    16'd9328: out <= 16'h0921;    16'd9329: out <= 16'h0386;    16'd9330: out <= 16'h05E2;    16'd9331: out <= 16'h02A0;
    16'd9332: out <= 16'h0241;    16'd9333: out <= 16'h0A36;    16'd9334: out <= 16'h01EE;    16'd9335: out <= 16'h0130;
    16'd9336: out <= 16'h04C0;    16'd9337: out <= 16'h0BB7;    16'd9338: out <= 16'h054D;    16'd9339: out <= 16'hFBB8;
    16'd9340: out <= 16'h03A9;    16'd9341: out <= 16'h099E;    16'd9342: out <= 16'h0141;    16'd9343: out <= 16'h05D8;
    16'd9344: out <= 16'h00CE;    16'd9345: out <= 16'h0295;    16'd9346: out <= 16'h0EFF;    16'd9347: out <= 16'h05A9;
    16'd9348: out <= 16'h007C;    16'd9349: out <= 16'h0037;    16'd9350: out <= 16'h023B;    16'd9351: out <= 16'h0250;
    16'd9352: out <= 16'hFEB6;    16'd9353: out <= 16'h078A;    16'd9354: out <= 16'h0235;    16'd9355: out <= 16'h075A;
    16'd9356: out <= 16'h04AD;    16'd9357: out <= 16'h09A4;    16'd9358: out <= 16'hFD5E;    16'd9359: out <= 16'h0245;
    16'd9360: out <= 16'hFFF9;    16'd9361: out <= 16'h0432;    16'd9362: out <= 16'h0559;    16'd9363: out <= 16'h037A;
    16'd9364: out <= 16'h04F9;    16'd9365: out <= 16'h0567;    16'd9366: out <= 16'h0008;    16'd9367: out <= 16'h03D7;
    16'd9368: out <= 16'h047B;    16'd9369: out <= 16'h0244;    16'd9370: out <= 16'h00B5;    16'd9371: out <= 16'hFF80;
    16'd9372: out <= 16'hFD0C;    16'd9373: out <= 16'h07E8;    16'd9374: out <= 16'h054C;    16'd9375: out <= 16'hFF56;
    16'd9376: out <= 16'h042C;    16'd9377: out <= 16'h004F;    16'd9378: out <= 16'h0456;    16'd9379: out <= 16'h0424;
    16'd9380: out <= 16'h04C4;    16'd9381: out <= 16'hFF46;    16'd9382: out <= 16'h0318;    16'd9383: out <= 16'hFEE0;
    16'd9384: out <= 16'h026A;    16'd9385: out <= 16'hFB35;    16'd9386: out <= 16'h02D9;    16'd9387: out <= 16'hFBF8;
    16'd9388: out <= 16'h062F;    16'd9389: out <= 16'h075E;    16'd9390: out <= 16'h0415;    16'd9391: out <= 16'h0875;
    16'd9392: out <= 16'h0577;    16'd9393: out <= 16'h04DF;    16'd9394: out <= 16'h0BDA;    16'd9395: out <= 16'h0630;
    16'd9396: out <= 16'hFF0E;    16'd9397: out <= 16'hFE23;    16'd9398: out <= 16'h01D6;    16'd9399: out <= 16'h0275;
    16'd9400: out <= 16'h04FC;    16'd9401: out <= 16'h0090;    16'd9402: out <= 16'hFEF5;    16'd9403: out <= 16'hFBAB;
    16'd9404: out <= 16'h057A;    16'd9405: out <= 16'h0359;    16'd9406: out <= 16'h0487;    16'd9407: out <= 16'hFFA9;
    16'd9408: out <= 16'h073C;    16'd9409: out <= 16'h06CB;    16'd9410: out <= 16'h0533;    16'd9411: out <= 16'h008E;
    16'd9412: out <= 16'h0582;    16'd9413: out <= 16'hFEA0;    16'd9414: out <= 16'hFFEA;    16'd9415: out <= 16'h0891;
    16'd9416: out <= 16'hFEB3;    16'd9417: out <= 16'h06F6;    16'd9418: out <= 16'h03F3;    16'd9419: out <= 16'h0D40;
    16'd9420: out <= 16'h033D;    16'd9421: out <= 16'hFF2B;    16'd9422: out <= 16'hFC53;    16'd9423: out <= 16'h06C9;
    16'd9424: out <= 16'hFB36;    16'd9425: out <= 16'hFFFB;    16'd9426: out <= 16'hFB4A;    16'd9427: out <= 16'h035C;
    16'd9428: out <= 16'hFF11;    16'd9429: out <= 16'hFDC1;    16'd9430: out <= 16'h0187;    16'd9431: out <= 16'h04C2;
    16'd9432: out <= 16'hFCEE;    16'd9433: out <= 16'h0695;    16'd9434: out <= 16'h016B;    16'd9435: out <= 16'h01E2;
    16'd9436: out <= 16'hFFE9;    16'd9437: out <= 16'h0020;    16'd9438: out <= 16'h02A7;    16'd9439: out <= 16'h026D;
    16'd9440: out <= 16'hFD34;    16'd9441: out <= 16'h0944;    16'd9442: out <= 16'hFA50;    16'd9443: out <= 16'hFE39;
    16'd9444: out <= 16'h0207;    16'd9445: out <= 16'h0351;    16'd9446: out <= 16'hFE14;    16'd9447: out <= 16'hFDB5;
    16'd9448: out <= 16'h01CD;    16'd9449: out <= 16'hFBC7;    16'd9450: out <= 16'hFC2E;    16'd9451: out <= 16'h00E0;
    16'd9452: out <= 16'h0132;    16'd9453: out <= 16'hF9DC;    16'd9454: out <= 16'hFF40;    16'd9455: out <= 16'hFAC0;
    16'd9456: out <= 16'hFD0D;    16'd9457: out <= 16'hFFEA;    16'd9458: out <= 16'hF940;    16'd9459: out <= 16'h0051;
    16'd9460: out <= 16'hFEF0;    16'd9461: out <= 16'h0300;    16'd9462: out <= 16'h06FA;    16'd9463: out <= 16'hFFBB;
    16'd9464: out <= 16'hFD3D;    16'd9465: out <= 16'hFE4E;    16'd9466: out <= 16'h026A;    16'd9467: out <= 16'hFB8C;
    16'd9468: out <= 16'hFEF4;    16'd9469: out <= 16'h06B7;    16'd9470: out <= 16'h06E4;    16'd9471: out <= 16'h020A;
    16'd9472: out <= 16'h00FA;    16'd9473: out <= 16'h09FC;    16'd9474: out <= 16'h03CE;    16'd9475: out <= 16'hFF67;
    16'd9476: out <= 16'hFCD1;    16'd9477: out <= 16'hFA64;    16'd9478: out <= 16'hFED3;    16'd9479: out <= 16'hFF6F;
    16'd9480: out <= 16'h0142;    16'd9481: out <= 16'h0073;    16'd9482: out <= 16'hFE47;    16'd9483: out <= 16'hFBE4;
    16'd9484: out <= 16'hFCC5;    16'd9485: out <= 16'h023E;    16'd9486: out <= 16'h007F;    16'd9487: out <= 16'hFA0A;
    16'd9488: out <= 16'h0036;    16'd9489: out <= 16'h0093;    16'd9490: out <= 16'hFC34;    16'd9491: out <= 16'h004F;
    16'd9492: out <= 16'h006E;    16'd9493: out <= 16'h03B0;    16'd9494: out <= 16'hFC90;    16'd9495: out <= 16'h0352;
    16'd9496: out <= 16'h00BF;    16'd9497: out <= 16'h0097;    16'd9498: out <= 16'hFE6B;    16'd9499: out <= 16'hFBE2;
    16'd9500: out <= 16'h0131;    16'd9501: out <= 16'h0500;    16'd9502: out <= 16'hFADD;    16'd9503: out <= 16'hFD96;
    16'd9504: out <= 16'h02F5;    16'd9505: out <= 16'hFAC8;    16'd9506: out <= 16'h044F;    16'd9507: out <= 16'h0655;
    16'd9508: out <= 16'h021C;    16'd9509: out <= 16'h066D;    16'd9510: out <= 16'hF61E;    16'd9511: out <= 16'h0599;
    16'd9512: out <= 16'h03DD;    16'd9513: out <= 16'h0484;    16'd9514: out <= 16'hFDB7;    16'd9515: out <= 16'hFEB2;
    16'd9516: out <= 16'h00FA;    16'd9517: out <= 16'h0362;    16'd9518: out <= 16'h04B4;    16'd9519: out <= 16'h0261;
    16'd9520: out <= 16'h079A;    16'd9521: out <= 16'h0634;    16'd9522: out <= 16'h010D;    16'd9523: out <= 16'h08E0;
    16'd9524: out <= 16'h067A;    16'd9525: out <= 16'h039E;    16'd9526: out <= 16'h04D2;    16'd9527: out <= 16'h0307;
    16'd9528: out <= 16'h0575;    16'd9529: out <= 16'h032D;    16'd9530: out <= 16'h02C0;    16'd9531: out <= 16'hFF57;
    16'd9532: out <= 16'h0400;    16'd9533: out <= 16'hFFA4;    16'd9534: out <= 16'h0504;    16'd9535: out <= 16'h0566;
    16'd9536: out <= 16'h061B;    16'd9537: out <= 16'h0074;    16'd9538: out <= 16'h05D4;    16'd9539: out <= 16'hFD27;
    16'd9540: out <= 16'h03A7;    16'd9541: out <= 16'h047C;    16'd9542: out <= 16'h0181;    16'd9543: out <= 16'h0940;
    16'd9544: out <= 16'h03F3;    16'd9545: out <= 16'hFE30;    16'd9546: out <= 16'h0969;    16'd9547: out <= 16'hF987;
    16'd9548: out <= 16'h0538;    16'd9549: out <= 16'h04BF;    16'd9550: out <= 16'h0397;    16'd9551: out <= 16'h03DB;
    16'd9552: out <= 16'h05E1;    16'd9553: out <= 16'h019F;    16'd9554: out <= 16'hFE93;    16'd9555: out <= 16'h0140;
    16'd9556: out <= 16'h07EB;    16'd9557: out <= 16'h01C6;    16'd9558: out <= 16'h0378;    16'd9559: out <= 16'h0403;
    16'd9560: out <= 16'h065A;    16'd9561: out <= 16'h0808;    16'd9562: out <= 16'h0258;    16'd9563: out <= 16'h030E;
    16'd9564: out <= 16'h017D;    16'd9565: out <= 16'h04E1;    16'd9566: out <= 16'h0891;    16'd9567: out <= 16'h05EF;
    16'd9568: out <= 16'h0A45;    16'd9569: out <= 16'h0035;    16'd9570: out <= 16'h0438;    16'd9571: out <= 16'h03F3;
    16'd9572: out <= 16'h00C9;    16'd9573: out <= 16'h073F;    16'd9574: out <= 16'h05C6;    16'd9575: out <= 16'h087C;
    16'd9576: out <= 16'hFFB3;    16'd9577: out <= 16'h01E9;    16'd9578: out <= 16'h059E;    16'd9579: out <= 16'h04D3;
    16'd9580: out <= 16'h0F4A;    16'd9581: out <= 16'hFF73;    16'd9582: out <= 16'h0070;    16'd9583: out <= 16'hFF69;
    16'd9584: out <= 16'h00A2;    16'd9585: out <= 16'h03C6;    16'd9586: out <= 16'h0121;    16'd9587: out <= 16'h077A;
    16'd9588: out <= 16'hFD29;    16'd9589: out <= 16'h02DB;    16'd9590: out <= 16'h081B;    16'd9591: out <= 16'h029A;
    16'd9592: out <= 16'h07F1;    16'd9593: out <= 16'h05FE;    16'd9594: out <= 16'h018F;    16'd9595: out <= 16'h0236;
    16'd9596: out <= 16'hFD32;    16'd9597: out <= 16'h030B;    16'd9598: out <= 16'h081E;    16'd9599: out <= 16'h0AA6;
    16'd9600: out <= 16'h0472;    16'd9601: out <= 16'h07E7;    16'd9602: out <= 16'h04E3;    16'd9603: out <= 16'hFF80;
    16'd9604: out <= 16'h0674;    16'd9605: out <= 16'h0962;    16'd9606: out <= 16'h0537;    16'd9607: out <= 16'h08AD;
    16'd9608: out <= 16'h0460;    16'd9609: out <= 16'h0956;    16'd9610: out <= 16'h062E;    16'd9611: out <= 16'h073B;
    16'd9612: out <= 16'h0601;    16'd9613: out <= 16'h0632;    16'd9614: out <= 16'h03FF;    16'd9615: out <= 16'h01E4;
    16'd9616: out <= 16'h0327;    16'd9617: out <= 16'hFD8B;    16'd9618: out <= 16'h0067;    16'd9619: out <= 16'h06ED;
    16'd9620: out <= 16'h022A;    16'd9621: out <= 16'h0242;    16'd9622: out <= 16'h01FB;    16'd9623: out <= 16'h039C;
    16'd9624: out <= 16'h05BC;    16'd9625: out <= 16'h0063;    16'd9626: out <= 16'h07ED;    16'd9627: out <= 16'hF5EA;
    16'd9628: out <= 16'h075F;    16'd9629: out <= 16'h067D;    16'd9630: out <= 16'h00D5;    16'd9631: out <= 16'h096D;
    16'd9632: out <= 16'h0185;    16'd9633: out <= 16'h0886;    16'd9634: out <= 16'h019B;    16'd9635: out <= 16'h0652;
    16'd9636: out <= 16'h03F4;    16'd9637: out <= 16'h0907;    16'd9638: out <= 16'h055A;    16'd9639: out <= 16'hFF86;
    16'd9640: out <= 16'h0274;    16'd9641: out <= 16'h0459;    16'd9642: out <= 16'h0767;    16'd9643: out <= 16'hFF5F;
    16'd9644: out <= 16'h0482;    16'd9645: out <= 16'h00C2;    16'd9646: out <= 16'hFF8C;    16'd9647: out <= 16'h0A43;
    16'd9648: out <= 16'h07EF;    16'd9649: out <= 16'h0881;    16'd9650: out <= 16'h0086;    16'd9651: out <= 16'h03A6;
    16'd9652: out <= 16'h0327;    16'd9653: out <= 16'hFAA5;    16'd9654: out <= 16'h064F;    16'd9655: out <= 16'h028E;
    16'd9656: out <= 16'h056D;    16'd9657: out <= 16'h05CA;    16'd9658: out <= 16'h0868;    16'd9659: out <= 16'h0260;
    16'd9660: out <= 16'h052A;    16'd9661: out <= 16'h04E5;    16'd9662: out <= 16'h06D9;    16'd9663: out <= 16'h0ADF;
    16'd9664: out <= 16'h01E8;    16'd9665: out <= 16'h09FB;    16'd9666: out <= 16'h0126;    16'd9667: out <= 16'h099C;
    16'd9668: out <= 16'h0052;    16'd9669: out <= 16'hFC6D;    16'd9670: out <= 16'h0657;    16'd9671: out <= 16'h09B7;
    16'd9672: out <= 16'h025F;    16'd9673: out <= 16'h061F;    16'd9674: out <= 16'h034C;    16'd9675: out <= 16'h0E0F;
    16'd9676: out <= 16'h0162;    16'd9677: out <= 16'hFEBA;    16'd9678: out <= 16'hFEE5;    16'd9679: out <= 16'hFE11;
    16'd9680: out <= 16'hFBD2;    16'd9681: out <= 16'h01FD;    16'd9682: out <= 16'hFB06;    16'd9683: out <= 16'h0284;
    16'd9684: out <= 16'hFE1B;    16'd9685: out <= 16'h04A0;    16'd9686: out <= 16'hFF51;    16'd9687: out <= 16'hFE5C;
    16'd9688: out <= 16'hFEAF;    16'd9689: out <= 16'h018C;    16'd9690: out <= 16'h016A;    16'd9691: out <= 16'h002E;
    16'd9692: out <= 16'hFDE4;    16'd9693: out <= 16'h01AF;    16'd9694: out <= 16'h03D4;    16'd9695: out <= 16'h050D;
    16'd9696: out <= 16'hFDCD;    16'd9697: out <= 16'hFB86;    16'd9698: out <= 16'h05FD;    16'd9699: out <= 16'h036C;
    16'd9700: out <= 16'hFD00;    16'd9701: out <= 16'h013C;    16'd9702: out <= 16'h043D;    16'd9703: out <= 16'h0172;
    16'd9704: out <= 16'h01FC;    16'd9705: out <= 16'h0154;    16'd9706: out <= 16'h0403;    16'd9707: out <= 16'hF75B;
    16'd9708: out <= 16'h0254;    16'd9709: out <= 16'hF953;    16'd9710: out <= 16'h00F2;    16'd9711: out <= 16'h03CB;
    16'd9712: out <= 16'hFED8;    16'd9713: out <= 16'h058B;    16'd9714: out <= 16'hFB89;    16'd9715: out <= 16'hFF0F;
    16'd9716: out <= 16'h0359;    16'd9717: out <= 16'hFD15;    16'd9718: out <= 16'h0358;    16'd9719: out <= 16'hFEF3;
    16'd9720: out <= 16'h005E;    16'd9721: out <= 16'hFFAA;    16'd9722: out <= 16'hF99A;    16'd9723: out <= 16'h0432;
    16'd9724: out <= 16'hFB4D;    16'd9725: out <= 16'hFCA1;    16'd9726: out <= 16'hFF0A;    16'd9727: out <= 16'h05C0;
    16'd9728: out <= 16'hFB54;    16'd9729: out <= 16'h01A5;    16'd9730: out <= 16'h0066;    16'd9731: out <= 16'h0126;
    16'd9732: out <= 16'hFBE4;    16'd9733: out <= 16'h027F;    16'd9734: out <= 16'hFB95;    16'd9735: out <= 16'h0282;
    16'd9736: out <= 16'h0739;    16'd9737: out <= 16'h0198;    16'd9738: out <= 16'h0A76;    16'd9739: out <= 16'h0175;
    16'd9740: out <= 16'h04C7;    16'd9741: out <= 16'hF88B;    16'd9742: out <= 16'hFC38;    16'd9743: out <= 16'h0239;
    16'd9744: out <= 16'hFF83;    16'd9745: out <= 16'h0047;    16'd9746: out <= 16'hFD53;    16'd9747: out <= 16'h03F7;
    16'd9748: out <= 16'hF9DA;    16'd9749: out <= 16'h0310;    16'd9750: out <= 16'h0258;    16'd9751: out <= 16'hFF7E;
    16'd9752: out <= 16'h0001;    16'd9753: out <= 16'h033D;    16'd9754: out <= 16'h0089;    16'd9755: out <= 16'h0513;
    16'd9756: out <= 16'hF6CD;    16'd9757: out <= 16'h04D5;    16'd9758: out <= 16'h0062;    16'd9759: out <= 16'hFF39;
    16'd9760: out <= 16'hFC4C;    16'd9761: out <= 16'h05D7;    16'd9762: out <= 16'h00BF;    16'd9763: out <= 16'hFF11;
    16'd9764: out <= 16'h013A;    16'd9765: out <= 16'hFE7A;    16'd9766: out <= 16'hFBDE;    16'd9767: out <= 16'h074C;
    16'd9768: out <= 16'hFF93;    16'd9769: out <= 16'hFC6D;    16'd9770: out <= 16'h06F5;    16'd9771: out <= 16'h0000;
    16'd9772: out <= 16'h03B3;    16'd9773: out <= 16'h03D2;    16'd9774: out <= 16'h0079;    16'd9775: out <= 16'h0280;
    16'd9776: out <= 16'h019F;    16'd9777: out <= 16'hFDB2;    16'd9778: out <= 16'h0203;    16'd9779: out <= 16'h0256;
    16'd9780: out <= 16'h051E;    16'd9781: out <= 16'h0B18;    16'd9782: out <= 16'h03C8;    16'd9783: out <= 16'h0630;
    16'd9784: out <= 16'h0799;    16'd9785: out <= 16'hFBD9;    16'd9786: out <= 16'h055B;    16'd9787: out <= 16'h0D6C;
    16'd9788: out <= 16'h0211;    16'd9789: out <= 16'hFF65;    16'd9790: out <= 16'h0285;    16'd9791: out <= 16'h04B2;
    16'd9792: out <= 16'h09FF;    16'd9793: out <= 16'hFB7A;    16'd9794: out <= 16'h026B;    16'd9795: out <= 16'h04BC;
    16'd9796: out <= 16'h0B4B;    16'd9797: out <= 16'h04D6;    16'd9798: out <= 16'hFFD7;    16'd9799: out <= 16'h0136;
    16'd9800: out <= 16'h0592;    16'd9801: out <= 16'h052B;    16'd9802: out <= 16'h0297;    16'd9803: out <= 16'hFB6F;
    16'd9804: out <= 16'h0706;    16'd9805: out <= 16'hFC2E;    16'd9806: out <= 16'h0593;    16'd9807: out <= 16'h0326;
    16'd9808: out <= 16'h05FD;    16'd9809: out <= 16'h08ED;    16'd9810: out <= 16'h0423;    16'd9811: out <= 16'h048C;
    16'd9812: out <= 16'hFFEC;    16'd9813: out <= 16'h0609;    16'd9814: out <= 16'h0469;    16'd9815: out <= 16'h05CE;
    16'd9816: out <= 16'hFE12;    16'd9817: out <= 16'h021F;    16'd9818: out <= 16'h03CF;    16'd9819: out <= 16'hFFDB;
    16'd9820: out <= 16'h02E8;    16'd9821: out <= 16'h0515;    16'd9822: out <= 16'hFEEB;    16'd9823: out <= 16'h0587;
    16'd9824: out <= 16'h02A3;    16'd9825: out <= 16'h08DE;    16'd9826: out <= 16'h04E5;    16'd9827: out <= 16'hFD1E;
    16'd9828: out <= 16'hFCB2;    16'd9829: out <= 16'h0716;    16'd9830: out <= 16'h06EC;    16'd9831: out <= 16'hFFFB;
    16'd9832: out <= 16'hFDB1;    16'd9833: out <= 16'h05C1;    16'd9834: out <= 16'h06B2;    16'd9835: out <= 16'hFC9D;
    16'd9836: out <= 16'h02D3;    16'd9837: out <= 16'h0556;    16'd9838: out <= 16'h0520;    16'd9839: out <= 16'hFF95;
    16'd9840: out <= 16'h0557;    16'd9841: out <= 16'h07EE;    16'd9842: out <= 16'hFCC0;    16'd9843: out <= 16'h084F;
    16'd9844: out <= 16'h08DB;    16'd9845: out <= 16'h05F9;    16'd9846: out <= 16'h028C;    16'd9847: out <= 16'h06DF;
    16'd9848: out <= 16'h086F;    16'd9849: out <= 16'h058D;    16'd9850: out <= 16'h01C7;    16'd9851: out <= 16'h0141;
    16'd9852: out <= 16'hFF37;    16'd9853: out <= 16'h0261;    16'd9854: out <= 16'h0936;    16'd9855: out <= 16'h04E9;
    16'd9856: out <= 16'h0959;    16'd9857: out <= 16'h074B;    16'd9858: out <= 16'h0127;    16'd9859: out <= 16'h051A;
    16'd9860: out <= 16'hFFEC;    16'd9861: out <= 16'h0323;    16'd9862: out <= 16'h0405;    16'd9863: out <= 16'h0991;
    16'd9864: out <= 16'hFF11;    16'd9865: out <= 16'hFC91;    16'd9866: out <= 16'h03F2;    16'd9867: out <= 16'hFFF4;
    16'd9868: out <= 16'h0669;    16'd9869: out <= 16'h027D;    16'd9870: out <= 16'h067B;    16'd9871: out <= 16'h0760;
    16'd9872: out <= 16'h0835;    16'd9873: out <= 16'h061C;    16'd9874: out <= 16'h04CC;    16'd9875: out <= 16'h00F2;
    16'd9876: out <= 16'h01C2;    16'd9877: out <= 16'h0525;    16'd9878: out <= 16'h0631;    16'd9879: out <= 16'hFFCD;
    16'd9880: out <= 16'h01E1;    16'd9881: out <= 16'h0462;    16'd9882: out <= 16'h0148;    16'd9883: out <= 16'h03D0;
    16'd9884: out <= 16'h0A63;    16'd9885: out <= 16'h0861;    16'd9886: out <= 16'h05BB;    16'd9887: out <= 16'h03B8;
    16'd9888: out <= 16'h02FB;    16'd9889: out <= 16'hFE25;    16'd9890: out <= 16'h0775;    16'd9891: out <= 16'h053E;
    16'd9892: out <= 16'h0271;    16'd9893: out <= 16'h0767;    16'd9894: out <= 16'h022B;    16'd9895: out <= 16'h0470;
    16'd9896: out <= 16'h086D;    16'd9897: out <= 16'h05FC;    16'd9898: out <= 16'h0509;    16'd9899: out <= 16'h08CF;
    16'd9900: out <= 16'h04A3;    16'd9901: out <= 16'h0453;    16'd9902: out <= 16'h0641;    16'd9903: out <= 16'h0360;
    16'd9904: out <= 16'h03E6;    16'd9905: out <= 16'hFEF7;    16'd9906: out <= 16'h05F5;    16'd9907: out <= 16'h04BE;
    16'd9908: out <= 16'h02A3;    16'd9909: out <= 16'hFE86;    16'd9910: out <= 16'h0EFB;    16'd9911: out <= 16'h0472;
    16'd9912: out <= 16'h0B69;    16'd9913: out <= 16'hFD8A;    16'd9914: out <= 16'h00AC;    16'd9915: out <= 16'h023C;
    16'd9916: out <= 16'h06D9;    16'd9917: out <= 16'h0627;    16'd9918: out <= 16'h016B;    16'd9919: out <= 16'h05A9;
    16'd9920: out <= 16'hFF1A;    16'd9921: out <= 16'h088E;    16'd9922: out <= 16'h0A34;    16'd9923: out <= 16'h0560;
    16'd9924: out <= 16'h0412;    16'd9925: out <= 16'h0993;    16'd9926: out <= 16'h00AB;    16'd9927: out <= 16'h06C2;
    16'd9928: out <= 16'h01D7;    16'd9929: out <= 16'h0280;    16'd9930: out <= 16'hFA9A;    16'd9931: out <= 16'h020A;
    16'd9932: out <= 16'h0163;    16'd9933: out <= 16'h03D5;    16'd9934: out <= 16'h046B;    16'd9935: out <= 16'hFB6C;
    16'd9936: out <= 16'h0225;    16'd9937: out <= 16'h0203;    16'd9938: out <= 16'hFF45;    16'd9939: out <= 16'hFC6B;
    16'd9940: out <= 16'h014B;    16'd9941: out <= 16'h0018;    16'd9942: out <= 16'h016D;    16'd9943: out <= 16'h0322;
    16'd9944: out <= 16'hFF4D;    16'd9945: out <= 16'hFF15;    16'd9946: out <= 16'h09BF;    16'd9947: out <= 16'h0294;
    16'd9948: out <= 16'hFBE6;    16'd9949: out <= 16'h0306;    16'd9950: out <= 16'h057C;    16'd9951: out <= 16'hFCE3;
    16'd9952: out <= 16'hFCF1;    16'd9953: out <= 16'hFB46;    16'd9954: out <= 16'hFBDF;    16'd9955: out <= 16'hF914;
    16'd9956: out <= 16'hFE3E;    16'd9957: out <= 16'hFECE;    16'd9958: out <= 16'hFA96;    16'd9959: out <= 16'h0281;
    16'd9960: out <= 16'hFB02;    16'd9961: out <= 16'hF987;    16'd9962: out <= 16'h0215;    16'd9963: out <= 16'h029A;
    16'd9964: out <= 16'hFFC9;    16'd9965: out <= 16'hF2F2;    16'd9966: out <= 16'hFE59;    16'd9967: out <= 16'hFF90;
    16'd9968: out <= 16'h04CA;    16'd9969: out <= 16'h00BB;    16'd9970: out <= 16'h0246;    16'd9971: out <= 16'hFD80;
    16'd9972: out <= 16'hF8ED;    16'd9973: out <= 16'hFBE6;    16'd9974: out <= 16'hFD20;    16'd9975: out <= 16'hFDDB;
    16'd9976: out <= 16'h03F5;    16'd9977: out <= 16'h003B;    16'd9978: out <= 16'h058B;    16'd9979: out <= 16'h0156;
    16'd9980: out <= 16'h05EF;    16'd9981: out <= 16'hFBAE;    16'd9982: out <= 16'hFC6E;    16'd9983: out <= 16'h0129;
    16'd9984: out <= 16'h06E0;    16'd9985: out <= 16'hFECC;    16'd9986: out <= 16'hFFA4;    16'd9987: out <= 16'hF954;
    16'd9988: out <= 16'hFF75;    16'd9989: out <= 16'h00C3;    16'd9990: out <= 16'h02E6;    16'd9991: out <= 16'hFB12;
    16'd9992: out <= 16'h00B4;    16'd9993: out <= 16'h0651;    16'd9994: out <= 16'hFF05;    16'd9995: out <= 16'h00B0;
    16'd9996: out <= 16'hFD7D;    16'd9997: out <= 16'hFCCE;    16'd9998: out <= 16'hFDA7;    16'd9999: out <= 16'hFF27;
    16'd10000: out <= 16'h06B1;    16'd10001: out <= 16'h011F;    16'd10002: out <= 16'h0128;    16'd10003: out <= 16'h03D0;
    16'd10004: out <= 16'hFD6B;    16'd10005: out <= 16'h0086;    16'd10006: out <= 16'hFFB8;    16'd10007: out <= 16'h06E5;
    16'd10008: out <= 16'h01CC;    16'd10009: out <= 16'hFC1C;    16'd10010: out <= 16'hFDE9;    16'd10011: out <= 16'h04A5;
    16'd10012: out <= 16'h051A;    16'd10013: out <= 16'hFE3F;    16'd10014: out <= 16'h0437;    16'd10015: out <= 16'hFD60;
    16'd10016: out <= 16'h086D;    16'd10017: out <= 16'h0510;    16'd10018: out <= 16'hFD41;    16'd10019: out <= 16'hFBDA;
    16'd10020: out <= 16'hF534;    16'd10021: out <= 16'hFD7C;    16'd10022: out <= 16'h0226;    16'd10023: out <= 16'h010D;
    16'd10024: out <= 16'h0135;    16'd10025: out <= 16'hFD34;    16'd10026: out <= 16'h0257;    16'd10027: out <= 16'h034F;
    16'd10028: out <= 16'hFECD;    16'd10029: out <= 16'h01F9;    16'd10030: out <= 16'h05D8;    16'd10031: out <= 16'h03C3;
    16'd10032: out <= 16'h0299;    16'd10033: out <= 16'hFDE4;    16'd10034: out <= 16'h0303;    16'd10035: out <= 16'h0035;
    16'd10036: out <= 16'hFEAE;    16'd10037: out <= 16'h03F2;    16'd10038: out <= 16'h0367;    16'd10039: out <= 16'h048E;
    16'd10040: out <= 16'h0631;    16'd10041: out <= 16'h044F;    16'd10042: out <= 16'h04AA;    16'd10043: out <= 16'h0349;
    16'd10044: out <= 16'h01B8;    16'd10045: out <= 16'h05E5;    16'd10046: out <= 16'h0488;    16'd10047: out <= 16'h0580;
    16'd10048: out <= 16'h0054;    16'd10049: out <= 16'hF896;    16'd10050: out <= 16'h0264;    16'd10051: out <= 16'h0770;
    16'd10052: out <= 16'hFD4B;    16'd10053: out <= 16'h043D;    16'd10054: out <= 16'h0334;    16'd10055: out <= 16'h0934;
    16'd10056: out <= 16'h0309;    16'd10057: out <= 16'h0668;    16'd10058: out <= 16'h0722;    16'd10059: out <= 16'hFEA5;
    16'd10060: out <= 16'h003C;    16'd10061: out <= 16'h00A9;    16'd10062: out <= 16'h00CC;    16'd10063: out <= 16'hFF84;
    16'd10064: out <= 16'h04C2;    16'd10065: out <= 16'h00F9;    16'd10066: out <= 16'h044D;    16'd10067: out <= 16'h087F;
    16'd10068: out <= 16'h0251;    16'd10069: out <= 16'h0860;    16'd10070: out <= 16'h0B4F;    16'd10071: out <= 16'h010F;
    16'd10072: out <= 16'h05F6;    16'd10073: out <= 16'h0374;    16'd10074: out <= 16'h0292;    16'd10075: out <= 16'hFE70;
    16'd10076: out <= 16'h07D5;    16'd10077: out <= 16'h07AD;    16'd10078: out <= 16'h0048;    16'd10079: out <= 16'h0AD7;
    16'd10080: out <= 16'h054F;    16'd10081: out <= 16'h04C2;    16'd10082: out <= 16'h0354;    16'd10083: out <= 16'h0975;
    16'd10084: out <= 16'h011D;    16'd10085: out <= 16'h04C5;    16'd10086: out <= 16'h06E3;    16'd10087: out <= 16'h0369;
    16'd10088: out <= 16'h0565;    16'd10089: out <= 16'h060F;    16'd10090: out <= 16'h05E3;    16'd10091: out <= 16'h081B;
    16'd10092: out <= 16'h047E;    16'd10093: out <= 16'h02CD;    16'd10094: out <= 16'h0026;    16'd10095: out <= 16'h058B;
    16'd10096: out <= 16'h0455;    16'd10097: out <= 16'h081A;    16'd10098: out <= 16'h09C5;    16'd10099: out <= 16'h016E;
    16'd10100: out <= 16'h02BE;    16'd10101: out <= 16'h0923;    16'd10102: out <= 16'hFBD1;    16'd10103: out <= 16'h04C3;
    16'd10104: out <= 16'hFC80;    16'd10105: out <= 16'hFE8D;    16'd10106: out <= 16'h076B;    16'd10107: out <= 16'h04CB;
    16'd10108: out <= 16'hFFA8;    16'd10109: out <= 16'h0821;    16'd10110: out <= 16'h06A2;    16'd10111: out <= 16'h0D0A;
    16'd10112: out <= 16'h048E;    16'd10113: out <= 16'h037A;    16'd10114: out <= 16'hFCFC;    16'd10115: out <= 16'h0096;
    16'd10116: out <= 16'h03A0;    16'd10117: out <= 16'h0622;    16'd10118: out <= 16'h0264;    16'd10119: out <= 16'hFD85;
    16'd10120: out <= 16'h052B;    16'd10121: out <= 16'h05A6;    16'd10122: out <= 16'h0016;    16'd10123: out <= 16'h02B7;
    16'd10124: out <= 16'h0774;    16'd10125: out <= 16'h076F;    16'd10126: out <= 16'h01FF;    16'd10127: out <= 16'h03B1;
    16'd10128: out <= 16'hF93F;    16'd10129: out <= 16'hFFE4;    16'd10130: out <= 16'h08E6;    16'd10131: out <= 16'h0185;
    16'd10132: out <= 16'hF875;    16'd10133: out <= 16'h08DE;    16'd10134: out <= 16'h0510;    16'd10135: out <= 16'h099E;
    16'd10136: out <= 16'h075E;    16'd10137: out <= 16'h0367;    16'd10138: out <= 16'hFFBE;    16'd10139: out <= 16'h0B12;
    16'd10140: out <= 16'h0080;    16'd10141: out <= 16'h0601;    16'd10142: out <= 16'h062A;    16'd10143: out <= 16'hFBEC;
    16'd10144: out <= 16'h03A0;    16'd10145: out <= 16'hFB1C;    16'd10146: out <= 16'h0136;    16'd10147: out <= 16'h0635;
    16'd10148: out <= 16'h04C0;    16'd10149: out <= 16'h0BB6;    16'd10150: out <= 16'h074D;    16'd10151: out <= 16'h0792;
    16'd10152: out <= 16'hFEB0;    16'd10153: out <= 16'hFF0F;    16'd10154: out <= 16'h0102;    16'd10155: out <= 16'h02B1;
    16'd10156: out <= 16'h0886;    16'd10157: out <= 16'h016F;    16'd10158: out <= 16'h03B2;    16'd10159: out <= 16'hFD37;
    16'd10160: out <= 16'h049E;    16'd10161: out <= 16'h0255;    16'd10162: out <= 16'h0168;    16'd10163: out <= 16'h0440;
    16'd10164: out <= 16'hF8F1;    16'd10165: out <= 16'h024C;    16'd10166: out <= 16'h0351;    16'd10167: out <= 16'h04DE;
    16'd10168: out <= 16'h06AD;    16'd10169: out <= 16'h0C41;    16'd10170: out <= 16'h06E6;    16'd10171: out <= 16'h071D;
    16'd10172: out <= 16'hFF49;    16'd10173: out <= 16'h05EA;    16'd10174: out <= 16'h09E1;    16'd10175: out <= 16'h0274;
    16'd10176: out <= 16'h0257;    16'd10177: out <= 16'h06FF;    16'd10178: out <= 16'h04A7;    16'd10179: out <= 16'h05E7;
    16'd10180: out <= 16'hFD5D;    16'd10181: out <= 16'h0340;    16'd10182: out <= 16'h0049;    16'd10183: out <= 16'h0202;
    16'd10184: out <= 16'h0209;    16'd10185: out <= 16'h0870;    16'd10186: out <= 16'h04AF;    16'd10187: out <= 16'h0624;
    16'd10188: out <= 16'h0AB2;    16'd10189: out <= 16'h0122;    16'd10190: out <= 16'h0828;    16'd10191: out <= 16'h03A3;
    16'd10192: out <= 16'h0395;    16'd10193: out <= 16'h0483;    16'd10194: out <= 16'hFD19;    16'd10195: out <= 16'h0303;
    16'd10196: out <= 16'hFF35;    16'd10197: out <= 16'h05C1;    16'd10198: out <= 16'h000F;    16'd10199: out <= 16'hFD58;
    16'd10200: out <= 16'h03FB;    16'd10201: out <= 16'hFCF3;    16'd10202: out <= 16'hFC89;    16'd10203: out <= 16'hFD55;
    16'd10204: out <= 16'h02B7;    16'd10205: out <= 16'hFF8A;    16'd10206: out <= 16'h0269;    16'd10207: out <= 16'h02EA;
    16'd10208: out <= 16'hFD46;    16'd10209: out <= 16'h0081;    16'd10210: out <= 16'h0151;    16'd10211: out <= 16'hFE05;
    16'd10212: out <= 16'hFED8;    16'd10213: out <= 16'hFB7D;    16'd10214: out <= 16'hFFA4;    16'd10215: out <= 16'hFB55;
    16'd10216: out <= 16'hF9B6;    16'd10217: out <= 16'hFF94;    16'd10218: out <= 16'hFC6E;    16'd10219: out <= 16'h027A;
    16'd10220: out <= 16'h0324;    16'd10221: out <= 16'hFED5;    16'd10222: out <= 16'hFF9D;    16'd10223: out <= 16'hFFCB;
    16'd10224: out <= 16'h012D;    16'd10225: out <= 16'hFEDC;    16'd10226: out <= 16'h08F4;    16'd10227: out <= 16'h0603;
    16'd10228: out <= 16'h062C;    16'd10229: out <= 16'h0282;    16'd10230: out <= 16'h00D0;    16'd10231: out <= 16'hFC9D;
    16'd10232: out <= 16'h014D;    16'd10233: out <= 16'hFA82;    16'd10234: out <= 16'h00EF;    16'd10235: out <= 16'h0300;
    16'd10236: out <= 16'hF724;    16'd10237: out <= 16'h00E2;    16'd10238: out <= 16'hFCE0;    16'd10239: out <= 16'h0525;
    16'd10240: out <= 16'hFBE4;    16'd10241: out <= 16'hF825;    16'd10242: out <= 16'hFBEC;    16'd10243: out <= 16'h0520;
    16'd10244: out <= 16'hFD0D;    16'd10245: out <= 16'hFC8F;    16'd10246: out <= 16'hFAF2;    16'd10247: out <= 16'h014F;
    16'd10248: out <= 16'hFD6F;    16'd10249: out <= 16'h0A23;    16'd10250: out <= 16'h030A;    16'd10251: out <= 16'hF9CC;
    16'd10252: out <= 16'hFEC5;    16'd10253: out <= 16'hFEF2;    16'd10254: out <= 16'h00C5;    16'd10255: out <= 16'h0662;
    16'd10256: out <= 16'h006F;    16'd10257: out <= 16'h005E;    16'd10258: out <= 16'hFF54;    16'd10259: out <= 16'hFBA2;
    16'd10260: out <= 16'hFEA5;    16'd10261: out <= 16'hFDBF;    16'd10262: out <= 16'hF9B0;    16'd10263: out <= 16'hFA95;
    16'd10264: out <= 16'hFB76;    16'd10265: out <= 16'hF949;    16'd10266: out <= 16'h036F;    16'd10267: out <= 16'hFEEB;
    16'd10268: out <= 16'hFF02;    16'd10269: out <= 16'h02EF;    16'd10270: out <= 16'h0327;    16'd10271: out <= 16'h08CD;
    16'd10272: out <= 16'h0073;    16'd10273: out <= 16'hFB86;    16'd10274: out <= 16'h0373;    16'd10275: out <= 16'h0739;
    16'd10276: out <= 16'h00CC;    16'd10277: out <= 16'h070F;    16'd10278: out <= 16'h06A7;    16'd10279: out <= 16'hFC2D;
    16'd10280: out <= 16'hFA65;    16'd10281: out <= 16'hFD5C;    16'd10282: out <= 16'h045A;    16'd10283: out <= 16'h02D8;
    16'd10284: out <= 16'h0331;    16'd10285: out <= 16'h008C;    16'd10286: out <= 16'hFFB4;    16'd10287: out <= 16'h02E9;
    16'd10288: out <= 16'h0335;    16'd10289: out <= 16'h0C51;    16'd10290: out <= 16'hFD18;    16'd10291: out <= 16'h0860;
    16'd10292: out <= 16'h020D;    16'd10293: out <= 16'hFF07;    16'd10294: out <= 16'h0727;    16'd10295: out <= 16'h0813;
    16'd10296: out <= 16'h0970;    16'd10297: out <= 16'h07D4;    16'd10298: out <= 16'h07AF;    16'd10299: out <= 16'h0382;
    16'd10300: out <= 16'h0C12;    16'd10301: out <= 16'h0917;    16'd10302: out <= 16'h022D;    16'd10303: out <= 16'h00B1;
    16'd10304: out <= 16'h063E;    16'd10305: out <= 16'h04CF;    16'd10306: out <= 16'h02E1;    16'd10307: out <= 16'hFD01;
    16'd10308: out <= 16'h01DC;    16'd10309: out <= 16'h0863;    16'd10310: out <= 16'h0761;    16'd10311: out <= 16'h0231;
    16'd10312: out <= 16'h0532;    16'd10313: out <= 16'hFD8E;    16'd10314: out <= 16'h0204;    16'd10315: out <= 16'h054E;
    16'd10316: out <= 16'h046C;    16'd10317: out <= 16'hFDC5;    16'd10318: out <= 16'hFFD7;    16'd10319: out <= 16'h09F8;
    16'd10320: out <= 16'h0B2F;    16'd10321: out <= 16'hFBB7;    16'd10322: out <= 16'h038C;    16'd10323: out <= 16'h0585;
    16'd10324: out <= 16'h02C4;    16'd10325: out <= 16'h0179;    16'd10326: out <= 16'hFEB8;    16'd10327: out <= 16'h0770;
    16'd10328: out <= 16'h0146;    16'd10329: out <= 16'h00FA;    16'd10330: out <= 16'h01A8;    16'd10331: out <= 16'h029A;
    16'd10332: out <= 16'h04E3;    16'd10333: out <= 16'hFA8C;    16'd10334: out <= 16'h016B;    16'd10335: out <= 16'hFFA7;
    16'd10336: out <= 16'h0088;    16'd10337: out <= 16'hFF8D;    16'd10338: out <= 16'h000C;    16'd10339: out <= 16'h06D2;
    16'd10340: out <= 16'h005F;    16'd10341: out <= 16'h044C;    16'd10342: out <= 16'h0509;    16'd10343: out <= 16'h00C1;
    16'd10344: out <= 16'h04E5;    16'd10345: out <= 16'h07B1;    16'd10346: out <= 16'hFCF6;    16'd10347: out <= 16'h08CB;
    16'd10348: out <= 16'hFCA3;    16'd10349: out <= 16'h0765;    16'd10350: out <= 16'h01B5;    16'd10351: out <= 16'h00F0;
    16'd10352: out <= 16'hFFA3;    16'd10353: out <= 16'h043F;    16'd10354: out <= 16'h01FB;    16'd10355: out <= 16'hFCE4;
    16'd10356: out <= 16'hFF46;    16'd10357: out <= 16'h058D;    16'd10358: out <= 16'hFFBF;    16'd10359: out <= 16'h03C0;
    16'd10360: out <= 16'h03FD;    16'd10361: out <= 16'h0729;    16'd10362: out <= 16'h06F5;    16'd10363: out <= 16'h01FB;
    16'd10364: out <= 16'h051A;    16'd10365: out <= 16'h062C;    16'd10366: out <= 16'h04B2;    16'd10367: out <= 16'hFCD3;
    16'd10368: out <= 16'h01DF;    16'd10369: out <= 16'h0605;    16'd10370: out <= 16'h00A3;    16'd10371: out <= 16'h01C2;
    16'd10372: out <= 16'h074F;    16'd10373: out <= 16'h09E5;    16'd10374: out <= 16'h04DB;    16'd10375: out <= 16'h0251;
    16'd10376: out <= 16'h019A;    16'd10377: out <= 16'h034A;    16'd10378: out <= 16'h0445;    16'd10379: out <= 16'h0A94;
    16'd10380: out <= 16'h0561;    16'd10381: out <= 16'h0669;    16'd10382: out <= 16'h0289;    16'd10383: out <= 16'h0A16;
    16'd10384: out <= 16'hF8E5;    16'd10385: out <= 16'h09E2;    16'd10386: out <= 16'hFFF9;    16'd10387: out <= 16'h0426;
    16'd10388: out <= 16'h014D;    16'd10389: out <= 16'h0144;    16'd10390: out <= 16'h0860;    16'd10391: out <= 16'h023B;
    16'd10392: out <= 16'h09E1;    16'd10393: out <= 16'h0183;    16'd10394: out <= 16'h0BA5;    16'd10395: out <= 16'h05FE;
    16'd10396: out <= 16'h0908;    16'd10397: out <= 16'h00E6;    16'd10398: out <= 16'h0342;    16'd10399: out <= 16'h037D;
    16'd10400: out <= 16'h0136;    16'd10401: out <= 16'hFA21;    16'd10402: out <= 16'hFFE8;    16'd10403: out <= 16'h039C;
    16'd10404: out <= 16'h0097;    16'd10405: out <= 16'h029C;    16'd10406: out <= 16'h0378;    16'd10407: out <= 16'h0A17;
    16'd10408: out <= 16'h096B;    16'd10409: out <= 16'h0A20;    16'd10410: out <= 16'h0472;    16'd10411: out <= 16'hFE41;
    16'd10412: out <= 16'hFFD0;    16'd10413: out <= 16'h05DF;    16'd10414: out <= 16'h019F;    16'd10415: out <= 16'h01CB;
    16'd10416: out <= 16'h020B;    16'd10417: out <= 16'h0345;    16'd10418: out <= 16'h0087;    16'd10419: out <= 16'h06DC;
    16'd10420: out <= 16'h02AB;    16'd10421: out <= 16'h0704;    16'd10422: out <= 16'h01FF;    16'd10423: out <= 16'h0431;
    16'd10424: out <= 16'h0676;    16'd10425: out <= 16'h08D9;    16'd10426: out <= 16'h082F;    16'd10427: out <= 16'hFF13;
    16'd10428: out <= 16'h0960;    16'd10429: out <= 16'hFE9A;    16'd10430: out <= 16'h00F1;    16'd10431: out <= 16'hFF8F;
    16'd10432: out <= 16'h00B5;    16'd10433: out <= 16'h05C6;    16'd10434: out <= 16'h06A8;    16'd10435: out <= 16'h05CA;
    16'd10436: out <= 16'h0333;    16'd10437: out <= 16'hFF19;    16'd10438: out <= 16'h0222;    16'd10439: out <= 16'h03DD;
    16'd10440: out <= 16'h0563;    16'd10441: out <= 16'h0336;    16'd10442: out <= 16'h044F;    16'd10443: out <= 16'h01DA;
    16'd10444: out <= 16'h074F;    16'd10445: out <= 16'h0AB8;    16'd10446: out <= 16'h0089;    16'd10447: out <= 16'h01E8;
    16'd10448: out <= 16'h038C;    16'd10449: out <= 16'hFE70;    16'd10450: out <= 16'h020A;    16'd10451: out <= 16'h0371;
    16'd10452: out <= 16'hFCB6;    16'd10453: out <= 16'h001E;    16'd10454: out <= 16'h0319;    16'd10455: out <= 16'hFBAA;
    16'd10456: out <= 16'hFC6F;    16'd10457: out <= 16'hFBE7;    16'd10458: out <= 16'hFA0A;    16'd10459: out <= 16'h00E5;
    16'd10460: out <= 16'hFC58;    16'd10461: out <= 16'hFBA6;    16'd10462: out <= 16'hFC98;    16'd10463: out <= 16'hF6B8;
    16'd10464: out <= 16'hFDEA;    16'd10465: out <= 16'h027E;    16'd10466: out <= 16'h0075;    16'd10467: out <= 16'hFD97;
    16'd10468: out <= 16'h0245;    16'd10469: out <= 16'hFEDF;    16'd10470: out <= 16'h028B;    16'd10471: out <= 16'h0205;
    16'd10472: out <= 16'h041F;    16'd10473: out <= 16'hFED0;    16'd10474: out <= 16'h046B;    16'd10475: out <= 16'hFB6A;
    16'd10476: out <= 16'hFC97;    16'd10477: out <= 16'hFC46;    16'd10478: out <= 16'hFEEA;    16'd10479: out <= 16'h07B4;
    16'd10480: out <= 16'h0185;    16'd10481: out <= 16'hFD9A;    16'd10482: out <= 16'hFF97;    16'd10483: out <= 16'hFCDB;
    16'd10484: out <= 16'h0030;    16'd10485: out <= 16'hFAF6;    16'd10486: out <= 16'hFD05;    16'd10487: out <= 16'h024B;
    16'd10488: out <= 16'hFD5C;    16'd10489: out <= 16'h00C3;    16'd10490: out <= 16'hFE28;    16'd10491: out <= 16'hFCC5;
    16'd10492: out <= 16'h08BB;    16'd10493: out <= 16'h01B9;    16'd10494: out <= 16'h05B9;    16'd10495: out <= 16'h0244;
    16'd10496: out <= 16'hFE82;    16'd10497: out <= 16'hFF63;    16'd10498: out <= 16'h0056;    16'd10499: out <= 16'h072A;
    16'd10500: out <= 16'hFE10;    16'd10501: out <= 16'h0237;    16'd10502: out <= 16'h0254;    16'd10503: out <= 16'h01A8;
    16'd10504: out <= 16'hFEE1;    16'd10505: out <= 16'hF809;    16'd10506: out <= 16'hF91D;    16'd10507: out <= 16'h016C;
    16'd10508: out <= 16'hFBD3;    16'd10509: out <= 16'h018C;    16'd10510: out <= 16'hFEFC;    16'd10511: out <= 16'h045E;
    16'd10512: out <= 16'hFF9C;    16'd10513: out <= 16'h0322;    16'd10514: out <= 16'h051E;    16'd10515: out <= 16'h0123;
    16'd10516: out <= 16'hFD3B;    16'd10517: out <= 16'h049E;    16'd10518: out <= 16'hFEDE;    16'd10519: out <= 16'h048E;
    16'd10520: out <= 16'hFAA3;    16'd10521: out <= 16'hFAF1;    16'd10522: out <= 16'h0034;    16'd10523: out <= 16'hFA98;
    16'd10524: out <= 16'h03B6;    16'd10525: out <= 16'h077A;    16'd10526: out <= 16'hFA25;    16'd10527: out <= 16'h004C;
    16'd10528: out <= 16'hFF39;    16'd10529: out <= 16'hFEF6;    16'd10530: out <= 16'hF734;    16'd10531: out <= 16'hFCF1;
    16'd10532: out <= 16'hFEED;    16'd10533: out <= 16'h05A3;    16'd10534: out <= 16'h0913;    16'd10535: out <= 16'hFF22;
    16'd10536: out <= 16'h02B4;    16'd10537: out <= 16'h0241;    16'd10538: out <= 16'h089A;    16'd10539: out <= 16'h00C0;
    16'd10540: out <= 16'h0621;    16'd10541: out <= 16'h0628;    16'd10542: out <= 16'h0B1C;    16'd10543: out <= 16'h0245;
    16'd10544: out <= 16'h02F8;    16'd10545: out <= 16'h0078;    16'd10546: out <= 16'h011F;    16'd10547: out <= 16'h07F7;
    16'd10548: out <= 16'h0378;    16'd10549: out <= 16'h075A;    16'd10550: out <= 16'h0751;    16'd10551: out <= 16'h009C;
    16'd10552: out <= 16'h0211;    16'd10553: out <= 16'h05E1;    16'd10554: out <= 16'hF993;    16'd10555: out <= 16'hFB1D;
    16'd10556: out <= 16'h01E9;    16'd10557: out <= 16'h02DC;    16'd10558: out <= 16'h0344;    16'd10559: out <= 16'h0580;
    16'd10560: out <= 16'h021F;    16'd10561: out <= 16'h051A;    16'd10562: out <= 16'h06F9;    16'd10563: out <= 16'h07CA;
    16'd10564: out <= 16'h06FF;    16'd10565: out <= 16'hFF25;    16'd10566: out <= 16'h0781;    16'd10567: out <= 16'h05EF;
    16'd10568: out <= 16'h008F;    16'd10569: out <= 16'h0385;    16'd10570: out <= 16'h0080;    16'd10571: out <= 16'h0F96;
    16'd10572: out <= 16'h03C0;    16'd10573: out <= 16'h01DE;    16'd10574: out <= 16'hFF07;    16'd10575: out <= 16'hFD82;
    16'd10576: out <= 16'hFA89;    16'd10577: out <= 16'h012F;    16'd10578: out <= 16'h00D9;    16'd10579: out <= 16'h044E;
    16'd10580: out <= 16'h0D4C;    16'd10581: out <= 16'hFEE4;    16'd10582: out <= 16'h039A;    16'd10583: out <= 16'h0083;
    16'd10584: out <= 16'hFF97;    16'd10585: out <= 16'h0641;    16'd10586: out <= 16'h021B;    16'd10587: out <= 16'h02D2;
    16'd10588: out <= 16'h0384;    16'd10589: out <= 16'h0C9E;    16'd10590: out <= 16'h01CD;    16'd10591: out <= 16'h0134;
    16'd10592: out <= 16'h0A4E;    16'd10593: out <= 16'h07BA;    16'd10594: out <= 16'h0097;    16'd10595: out <= 16'h0378;
    16'd10596: out <= 16'h0792;    16'd10597: out <= 16'h03C0;    16'd10598: out <= 16'h0342;    16'd10599: out <= 16'hFC46;
    16'd10600: out <= 16'h045A;    16'd10601: out <= 16'h03A7;    16'd10602: out <= 16'h042C;    16'd10603: out <= 16'h0433;
    16'd10604: out <= 16'h0857;    16'd10605: out <= 16'h083D;    16'd10606: out <= 16'h01B1;    16'd10607: out <= 16'h03BE;
    16'd10608: out <= 16'hFD16;    16'd10609: out <= 16'hFDEE;    16'd10610: out <= 16'hFD58;    16'd10611: out <= 16'h0C21;
    16'd10612: out <= 16'h01B8;    16'd10613: out <= 16'h00B7;    16'd10614: out <= 16'hFFB3;    16'd10615: out <= 16'h00E5;
    16'd10616: out <= 16'h062D;    16'd10617: out <= 16'h08E9;    16'd10618: out <= 16'h0A61;    16'd10619: out <= 16'h03C6;
    16'd10620: out <= 16'h051A;    16'd10621: out <= 16'h0003;    16'd10622: out <= 16'h099D;    16'd10623: out <= 16'h0073;
    16'd10624: out <= 16'h0752;    16'd10625: out <= 16'h06E1;    16'd10626: out <= 16'h009D;    16'd10627: out <= 16'h08D0;
    16'd10628: out <= 16'h0617;    16'd10629: out <= 16'h042F;    16'd10630: out <= 16'h041E;    16'd10631: out <= 16'h0098;
    16'd10632: out <= 16'h0395;    16'd10633: out <= 16'h03EA;    16'd10634: out <= 16'h0401;    16'd10635: out <= 16'h048B;
    16'd10636: out <= 16'h0622;    16'd10637: out <= 16'h080E;    16'd10638: out <= 16'h02D4;    16'd10639: out <= 16'h0295;
    16'd10640: out <= 16'h07C8;    16'd10641: out <= 16'hFEBC;    16'd10642: out <= 16'h032F;    16'd10643: out <= 16'h0467;
    16'd10644: out <= 16'h04D0;    16'd10645: out <= 16'h019B;    16'd10646: out <= 16'h09DA;    16'd10647: out <= 16'h0710;
    16'd10648: out <= 16'h03A9;    16'd10649: out <= 16'h06B5;    16'd10650: out <= 16'h0A05;    16'd10651: out <= 16'h0429;
    16'd10652: out <= 16'hFF73;    16'd10653: out <= 16'h06D3;    16'd10654: out <= 16'h0C3E;    16'd10655: out <= 16'hF9F3;
    16'd10656: out <= 16'h0299;    16'd10657: out <= 16'h00F7;    16'd10658: out <= 16'h01C2;    16'd10659: out <= 16'hFF58;
    16'd10660: out <= 16'hFF77;    16'd10661: out <= 16'h0176;    16'd10662: out <= 16'h047F;    16'd10663: out <= 16'h0416;
    16'd10664: out <= 16'h04FE;    16'd10665: out <= 16'hFF49;    16'd10666: out <= 16'h0850;    16'd10667: out <= 16'h02E1;
    16'd10668: out <= 16'hF972;    16'd10669: out <= 16'h031C;    16'd10670: out <= 16'h03B5;    16'd10671: out <= 16'h0250;
    16'd10672: out <= 16'hFE9B;    16'd10673: out <= 16'h0489;    16'd10674: out <= 16'h036E;    16'd10675: out <= 16'h02F1;
    16'd10676: out <= 16'hFDF2;    16'd10677: out <= 16'h04C1;    16'd10678: out <= 16'h0368;    16'd10679: out <= 16'hFF9C;
    16'd10680: out <= 16'h02D3;    16'd10681: out <= 16'h03CC;    16'd10682: out <= 16'h0366;    16'd10683: out <= 16'h0046;
    16'd10684: out <= 16'hFD55;    16'd10685: out <= 16'h0422;    16'd10686: out <= 16'h034F;    16'd10687: out <= 16'h0246;
    16'd10688: out <= 16'h036C;    16'd10689: out <= 16'h08EF;    16'd10690: out <= 16'h00F5;    16'd10691: out <= 16'h03C3;
    16'd10692: out <= 16'hFFEF;    16'd10693: out <= 16'h0699;    16'd10694: out <= 16'h058F;    16'd10695: out <= 16'h0496;
    16'd10696: out <= 16'h016B;    16'd10697: out <= 16'h038C;    16'd10698: out <= 16'h04F9;    16'd10699: out <= 16'h017B;
    16'd10700: out <= 16'h0A2B;    16'd10701: out <= 16'h0314;    16'd10702: out <= 16'h06B3;    16'd10703: out <= 16'h05A9;
    16'd10704: out <= 16'h0536;    16'd10705: out <= 16'h039F;    16'd10706: out <= 16'h0009;    16'd10707: out <= 16'hFCE6;
    16'd10708: out <= 16'h05AB;    16'd10709: out <= 16'hFBD6;    16'd10710: out <= 16'h05CB;    16'd10711: out <= 16'h013E;
    16'd10712: out <= 16'h047E;    16'd10713: out <= 16'h0090;    16'd10714: out <= 16'hFD7D;    16'd10715: out <= 16'h00AE;
    16'd10716: out <= 16'h011D;    16'd10717: out <= 16'hFC0D;    16'd10718: out <= 16'hFF4B;    16'd10719: out <= 16'h01E6;
    16'd10720: out <= 16'hFF49;    16'd10721: out <= 16'h023A;    16'd10722: out <= 16'h01E4;    16'd10723: out <= 16'hFF0A;
    16'd10724: out <= 16'h00F8;    16'd10725: out <= 16'hF947;    16'd10726: out <= 16'hFBCB;    16'd10727: out <= 16'hFBC1;
    16'd10728: out <= 16'h01A9;    16'd10729: out <= 16'hFD5F;    16'd10730: out <= 16'hFD70;    16'd10731: out <= 16'hFCCB;
    16'd10732: out <= 16'hFCF7;    16'd10733: out <= 16'h0A9F;    16'd10734: out <= 16'hFFDD;    16'd10735: out <= 16'hFFD3;
    16'd10736: out <= 16'hFEF7;    16'd10737: out <= 16'h0354;    16'd10738: out <= 16'h037B;    16'd10739: out <= 16'hFCF0;
    16'd10740: out <= 16'hFD9C;    16'd10741: out <= 16'hFFCC;    16'd10742: out <= 16'h0094;    16'd10743: out <= 16'hFF9A;
    16'd10744: out <= 16'h03B0;    16'd10745: out <= 16'hFC11;    16'd10746: out <= 16'h0000;    16'd10747: out <= 16'h03F1;
    16'd10748: out <= 16'hFE13;    16'd10749: out <= 16'h00CB;    16'd10750: out <= 16'hFEBA;    16'd10751: out <= 16'h0470;
    16'd10752: out <= 16'h0187;    16'd10753: out <= 16'h0669;    16'd10754: out <= 16'hFF01;    16'd10755: out <= 16'h026C;
    16'd10756: out <= 16'h0091;    16'd10757: out <= 16'hFF91;    16'd10758: out <= 16'h03FB;    16'd10759: out <= 16'h010A;
    16'd10760: out <= 16'hFC38;    16'd10761: out <= 16'h011F;    16'd10762: out <= 16'hFF21;    16'd10763: out <= 16'h03E6;
    16'd10764: out <= 16'h00B9;    16'd10765: out <= 16'h09C4;    16'd10766: out <= 16'hFD24;    16'd10767: out <= 16'hFDA8;
    16'd10768: out <= 16'hF88F;    16'd10769: out <= 16'h02B1;    16'd10770: out <= 16'hFF64;    16'd10771: out <= 16'hFD77;
    16'd10772: out <= 16'hFD71;    16'd10773: out <= 16'h0502;    16'd10774: out <= 16'hF79E;    16'd10775: out <= 16'h023A;
    16'd10776: out <= 16'h023F;    16'd10777: out <= 16'h059C;    16'd10778: out <= 16'h0104;    16'd10779: out <= 16'h03F7;
    16'd10780: out <= 16'h0193;    16'd10781: out <= 16'hFC13;    16'd10782: out <= 16'hFF4D;    16'd10783: out <= 16'hFB2A;
    16'd10784: out <= 16'hFE26;    16'd10785: out <= 16'h02B0;    16'd10786: out <= 16'h0434;    16'd10787: out <= 16'h0149;
    16'd10788: out <= 16'h039E;    16'd10789: out <= 16'h0629;    16'd10790: out <= 16'h0192;    16'd10791: out <= 16'h036E;
    16'd10792: out <= 16'hFA47;    16'd10793: out <= 16'hFFAE;    16'd10794: out <= 16'h0029;    16'd10795: out <= 16'h0663;
    16'd10796: out <= 16'h0891;    16'd10797: out <= 16'h005F;    16'd10798: out <= 16'h00B6;    16'd10799: out <= 16'h049E;
    16'd10800: out <= 16'h0414;    16'd10801: out <= 16'h06DE;    16'd10802: out <= 16'h0760;    16'd10803: out <= 16'h07AA;
    16'd10804: out <= 16'h06E8;    16'd10805: out <= 16'hFF93;    16'd10806: out <= 16'h0609;    16'd10807: out <= 16'h02A3;
    16'd10808: out <= 16'h0570;    16'd10809: out <= 16'hFDFD;    16'd10810: out <= 16'h0223;    16'd10811: out <= 16'h058B;
    16'd10812: out <= 16'h05A1;    16'd10813: out <= 16'h08C0;    16'd10814: out <= 16'h028B;    16'd10815: out <= 16'h0B31;
    16'd10816: out <= 16'hFEB8;    16'd10817: out <= 16'h02BB;    16'd10818: out <= 16'h0015;    16'd10819: out <= 16'h0A1E;
    16'd10820: out <= 16'hFE02;    16'd10821: out <= 16'h08EC;    16'd10822: out <= 16'hFE73;    16'd10823: out <= 16'h03C0;
    16'd10824: out <= 16'h0B19;    16'd10825: out <= 16'h0030;    16'd10826: out <= 16'h03BA;    16'd10827: out <= 16'h0387;
    16'd10828: out <= 16'h0088;    16'd10829: out <= 16'h05D5;    16'd10830: out <= 16'h073E;    16'd10831: out <= 16'h00E7;
    16'd10832: out <= 16'h0830;    16'd10833: out <= 16'h0108;    16'd10834: out <= 16'h07CC;    16'd10835: out <= 16'hFFE1;
    16'd10836: out <= 16'h056A;    16'd10837: out <= 16'hFF3A;    16'd10838: out <= 16'h0111;    16'd10839: out <= 16'h00B1;
    16'd10840: out <= 16'h0819;    16'd10841: out <= 16'h06C6;    16'd10842: out <= 16'h0549;    16'd10843: out <= 16'h08F6;
    16'd10844: out <= 16'h048F;    16'd10845: out <= 16'hFC0A;    16'd10846: out <= 16'h0964;    16'd10847: out <= 16'h0512;
    16'd10848: out <= 16'h0301;    16'd10849: out <= 16'hFED9;    16'd10850: out <= 16'h02B9;    16'd10851: out <= 16'h02C7;
    16'd10852: out <= 16'h01B4;    16'd10853: out <= 16'h017F;    16'd10854: out <= 16'h0349;    16'd10855: out <= 16'h054A;
    16'd10856: out <= 16'h085B;    16'd10857: out <= 16'hFEB4;    16'd10858: out <= 16'hFFB5;    16'd10859: out <= 16'hFBB1;
    16'd10860: out <= 16'h0531;    16'd10861: out <= 16'h08C9;    16'd10862: out <= 16'h053D;    16'd10863: out <= 16'h0501;
    16'd10864: out <= 16'h0AAF;    16'd10865: out <= 16'h042B;    16'd10866: out <= 16'h075D;    16'd10867: out <= 16'h0270;
    16'd10868: out <= 16'h00BA;    16'd10869: out <= 16'h067F;    16'd10870: out <= 16'hFEA3;    16'd10871: out <= 16'h0290;
    16'd10872: out <= 16'h086F;    16'd10873: out <= 16'h0BDB;    16'd10874: out <= 16'h03FA;    16'd10875: out <= 16'h0074;
    16'd10876: out <= 16'h0336;    16'd10877: out <= 16'h0111;    16'd10878: out <= 16'h02DF;    16'd10879: out <= 16'h035A;
    16'd10880: out <= 16'h0220;    16'd10881: out <= 16'h035E;    16'd10882: out <= 16'h037A;    16'd10883: out <= 16'h07B7;
    16'd10884: out <= 16'h0179;    16'd10885: out <= 16'h0257;    16'd10886: out <= 16'h0908;    16'd10887: out <= 16'h042F;
    16'd10888: out <= 16'h0026;    16'd10889: out <= 16'h022E;    16'd10890: out <= 16'h035E;    16'd10891: out <= 16'h0122;
    16'd10892: out <= 16'h08C3;    16'd10893: out <= 16'h0AE8;    16'd10894: out <= 16'h0113;    16'd10895: out <= 16'h06CD;
    16'd10896: out <= 16'h04D5;    16'd10897: out <= 16'hFFE0;    16'd10898: out <= 16'h071F;    16'd10899: out <= 16'h0AA6;
    16'd10900: out <= 16'h082C;    16'd10901: out <= 16'h0096;    16'd10902: out <= 16'h06CE;    16'd10903: out <= 16'h05EA;
    16'd10904: out <= 16'h0AC9;    16'd10905: out <= 16'hFC2F;    16'd10906: out <= 16'h069B;    16'd10907: out <= 16'h009C;
    16'd10908: out <= 16'h08CA;    16'd10909: out <= 16'h0A34;    16'd10910: out <= 16'h08A0;    16'd10911: out <= 16'h02F2;
    16'd10912: out <= 16'h0465;    16'd10913: out <= 16'h046B;    16'd10914: out <= 16'h0BD5;    16'd10915: out <= 16'hFFF3;
    16'd10916: out <= 16'hFA22;    16'd10917: out <= 16'h0157;    16'd10918: out <= 16'h002E;    16'd10919: out <= 16'hFED5;
    16'd10920: out <= 16'h0A25;    16'd10921: out <= 16'h03DD;    16'd10922: out <= 16'h043E;    16'd10923: out <= 16'h0106;
    16'd10924: out <= 16'h0A1F;    16'd10925: out <= 16'h0360;    16'd10926: out <= 16'h0959;    16'd10927: out <= 16'h044D;
    16'd10928: out <= 16'hFFF0;    16'd10929: out <= 16'h05F0;    16'd10930: out <= 16'h0803;    16'd10931: out <= 16'h022F;
    16'd10932: out <= 16'h072F;    16'd10933: out <= 16'h0279;    16'd10934: out <= 16'h069A;    16'd10935: out <= 16'h0481;
    16'd10936: out <= 16'h0795;    16'd10937: out <= 16'h020F;    16'd10938: out <= 16'h0731;    16'd10939: out <= 16'h0068;
    16'd10940: out <= 16'h0160;    16'd10941: out <= 16'hFEE4;    16'd10942: out <= 16'h0378;    16'd10943: out <= 16'h08DE;
    16'd10944: out <= 16'h022D;    16'd10945: out <= 16'h0480;    16'd10946: out <= 16'h0556;    16'd10947: out <= 16'hFE4C;
    16'd10948: out <= 16'h0721;    16'd10949: out <= 16'h0098;    16'd10950: out <= 16'h0786;    16'd10951: out <= 16'hFC34;
    16'd10952: out <= 16'h0964;    16'd10953: out <= 16'h0310;    16'd10954: out <= 16'h0367;    16'd10955: out <= 16'h06AD;
    16'd10956: out <= 16'h06D1;    16'd10957: out <= 16'h034E;    16'd10958: out <= 16'h05E1;    16'd10959: out <= 16'h0247;
    16'd10960: out <= 16'h03E8;    16'd10961: out <= 16'h0736;    16'd10962: out <= 16'hFF5F;    16'd10963: out <= 16'hFE71;
    16'd10964: out <= 16'hFEEB;    16'd10965: out <= 16'hFFA6;    16'd10966: out <= 16'hFCE4;    16'd10967: out <= 16'h0227;
    16'd10968: out <= 16'h02AD;    16'd10969: out <= 16'h01E4;    16'd10970: out <= 16'h0528;    16'd10971: out <= 16'h01A5;
    16'd10972: out <= 16'hF80F;    16'd10973: out <= 16'hFE79;    16'd10974: out <= 16'hFF3A;    16'd10975: out <= 16'hFE1C;
    16'd10976: out <= 16'hFDF1;    16'd10977: out <= 16'hFD16;    16'd10978: out <= 16'hFE2E;    16'd10979: out <= 16'h01F3;
    16'd10980: out <= 16'hFD29;    16'd10981: out <= 16'h034D;    16'd10982: out <= 16'hFFE8;    16'd10983: out <= 16'hFAF6;
    16'd10984: out <= 16'hFC40;    16'd10985: out <= 16'hFE89;    16'd10986: out <= 16'h079F;    16'd10987: out <= 16'hFD67;
    16'd10988: out <= 16'hFF5D;    16'd10989: out <= 16'h00E5;    16'd10990: out <= 16'hFA2B;    16'd10991: out <= 16'hFD93;
    16'd10992: out <= 16'hFE34;    16'd10993: out <= 16'hFE92;    16'd10994: out <= 16'h0027;    16'd10995: out <= 16'hF7EF;
    16'd10996: out <= 16'hFD65;    16'd10997: out <= 16'hFF47;    16'd10998: out <= 16'hFFB6;    16'd10999: out <= 16'h000C;
    16'd11000: out <= 16'h0147;    16'd11001: out <= 16'hFDCA;    16'd11002: out <= 16'h014D;    16'd11003: out <= 16'hFCF2;
    16'd11004: out <= 16'hFFAF;    16'd11005: out <= 16'h07B3;    16'd11006: out <= 16'h07A4;    16'd11007: out <= 16'hFEB6;
    16'd11008: out <= 16'hFFE8;    16'd11009: out <= 16'h03CE;    16'd11010: out <= 16'hFFCF;    16'd11011: out <= 16'hFDEA;
    16'd11012: out <= 16'h02C6;    16'd11013: out <= 16'h0182;    16'd11014: out <= 16'hF6AC;    16'd11015: out <= 16'h0319;
    16'd11016: out <= 16'h01F8;    16'd11017: out <= 16'hFF0D;    16'd11018: out <= 16'h00A0;    16'd11019: out <= 16'hFC7D;
    16'd11020: out <= 16'hFCA1;    16'd11021: out <= 16'hFBD5;    16'd11022: out <= 16'hFC05;    16'd11023: out <= 16'hFA8E;
    16'd11024: out <= 16'h004F;    16'd11025: out <= 16'h0212;    16'd11026: out <= 16'h0533;    16'd11027: out <= 16'hFE09;
    16'd11028: out <= 16'hFD35;    16'd11029: out <= 16'hFE1C;    16'd11030: out <= 16'h00F7;    16'd11031: out <= 16'h086F;
    16'd11032: out <= 16'h0145;    16'd11033: out <= 16'h03A4;    16'd11034: out <= 16'hFC24;    16'd11035: out <= 16'h0B00;
    16'd11036: out <= 16'hFDC3;    16'd11037: out <= 16'hFFE4;    16'd11038: out <= 16'hFBC0;    16'd11039: out <= 16'h0470;
    16'd11040: out <= 16'h002F;    16'd11041: out <= 16'h0286;    16'd11042: out <= 16'hFB36;    16'd11043: out <= 16'h03F4;
    16'd11044: out <= 16'h06A5;    16'd11045: out <= 16'hFF05;    16'd11046: out <= 16'hFDAF;    16'd11047: out <= 16'hFEC4;
    16'd11048: out <= 16'h0712;    16'd11049: out <= 16'h046A;    16'd11050: out <= 16'h0735;    16'd11051: out <= 16'h0BE2;
    16'd11052: out <= 16'h04BC;    16'd11053: out <= 16'h0271;    16'd11054: out <= 16'h0660;    16'd11055: out <= 16'h033E;
    16'd11056: out <= 16'h0958;    16'd11057: out <= 16'h00EF;    16'd11058: out <= 16'h06DD;    16'd11059: out <= 16'h0788;
    16'd11060: out <= 16'h0759;    16'd11061: out <= 16'h01C1;    16'd11062: out <= 16'h109C;    16'd11063: out <= 16'h0652;
    16'd11064: out <= 16'h0384;    16'd11065: out <= 16'h0375;    16'd11066: out <= 16'h04E2;    16'd11067: out <= 16'hFF00;
    16'd11068: out <= 16'h03C8;    16'd11069: out <= 16'h01D9;    16'd11070: out <= 16'h062B;    16'd11071: out <= 16'h0184;
    16'd11072: out <= 16'h049D;    16'd11073: out <= 16'h054C;    16'd11074: out <= 16'h0072;    16'd11075: out <= 16'hFCD4;
    16'd11076: out <= 16'h0611;    16'd11077: out <= 16'h06E6;    16'd11078: out <= 16'h00E6;    16'd11079: out <= 16'h079C;
    16'd11080: out <= 16'hFF0F;    16'd11081: out <= 16'h0502;    16'd11082: out <= 16'h0707;    16'd11083: out <= 16'h0363;
    16'd11084: out <= 16'h08D3;    16'd11085: out <= 16'h0DF4;    16'd11086: out <= 16'hFDB5;    16'd11087: out <= 16'hFEEC;
    16'd11088: out <= 16'h03DE;    16'd11089: out <= 16'h0583;    16'd11090: out <= 16'h017A;    16'd11091: out <= 16'h076D;
    16'd11092: out <= 16'h09C2;    16'd11093: out <= 16'h01C5;    16'd11094: out <= 16'h0368;    16'd11095: out <= 16'hF9EA;
    16'd11096: out <= 16'h0886;    16'd11097: out <= 16'h01A5;    16'd11098: out <= 16'h04C5;    16'd11099: out <= 16'h046C;
    16'd11100: out <= 16'h04BD;    16'd11101: out <= 16'h0A1B;    16'd11102: out <= 16'hFEEC;    16'd11103: out <= 16'h02C4;
    16'd11104: out <= 16'h008D;    16'd11105: out <= 16'h0776;    16'd11106: out <= 16'h055C;    16'd11107: out <= 16'h0658;
    16'd11108: out <= 16'h03CD;    16'd11109: out <= 16'h017A;    16'd11110: out <= 16'h03C9;    16'd11111: out <= 16'hFFF8;
    16'd11112: out <= 16'h0279;    16'd11113: out <= 16'h007D;    16'd11114: out <= 16'h0377;    16'd11115: out <= 16'h0075;
    16'd11116: out <= 16'h0AB8;    16'd11117: out <= 16'hFF81;    16'd11118: out <= 16'h0246;    16'd11119: out <= 16'h026C;
    16'd11120: out <= 16'h0563;    16'd11121: out <= 16'h085C;    16'd11122: out <= 16'h0664;    16'd11123: out <= 16'h03C2;
    16'd11124: out <= 16'h0515;    16'd11125: out <= 16'h0798;    16'd11126: out <= 16'hFC2C;    16'd11127: out <= 16'h0889;
    16'd11128: out <= 16'h063F;    16'd11129: out <= 16'h0029;    16'd11130: out <= 16'h0EED;    16'd11131: out <= 16'h0323;
    16'd11132: out <= 16'h01C7;    16'd11133: out <= 16'h0408;    16'd11134: out <= 16'h0AF2;    16'd11135: out <= 16'h0083;
    16'd11136: out <= 16'h02F6;    16'd11137: out <= 16'h0A3B;    16'd11138: out <= 16'h0D4B;    16'd11139: out <= 16'h0353;
    16'd11140: out <= 16'hFFAD;    16'd11141: out <= 16'h07F8;    16'd11142: out <= 16'hFBE8;    16'd11143: out <= 16'h05AE;
    16'd11144: out <= 16'h092E;    16'd11145: out <= 16'h0977;    16'd11146: out <= 16'h0808;    16'd11147: out <= 16'h0433;
    16'd11148: out <= 16'h067B;    16'd11149: out <= 16'h0200;    16'd11150: out <= 16'h03D0;    16'd11151: out <= 16'h05D4;
    16'd11152: out <= 16'h05DF;    16'd11153: out <= 16'hFFA4;    16'd11154: out <= 16'hF8C3;    16'd11155: out <= 16'hFFF0;
    16'd11156: out <= 16'h0291;    16'd11157: out <= 16'hFBEF;    16'd11158: out <= 16'h05E9;    16'd11159: out <= 16'h0607;
    16'd11160: out <= 16'h02D4;    16'd11161: out <= 16'h0466;    16'd11162: out <= 16'h06E4;    16'd11163: out <= 16'h07B1;
    16'd11164: out <= 16'h0435;    16'd11165: out <= 16'h01B7;    16'd11166: out <= 16'h0478;    16'd11167: out <= 16'h0170;
    16'd11168: out <= 16'h017F;    16'd11169: out <= 16'h0F6C;    16'd11170: out <= 16'h013A;    16'd11171: out <= 16'hFF31;
    16'd11172: out <= 16'h00E1;    16'd11173: out <= 16'h0360;    16'd11174: out <= 16'h0CE4;    16'd11175: out <= 16'hFB91;
    16'd11176: out <= 16'h0264;    16'd11177: out <= 16'h056D;    16'd11178: out <= 16'h0453;    16'd11179: out <= 16'h0408;
    16'd11180: out <= 16'h00EC;    16'd11181: out <= 16'hFEAA;    16'd11182: out <= 16'h04C0;    16'd11183: out <= 16'h03F9;
    16'd11184: out <= 16'h0C75;    16'd11185: out <= 16'h0280;    16'd11186: out <= 16'h036F;    16'd11187: out <= 16'h087B;
    16'd11188: out <= 16'h0BFF;    16'd11189: out <= 16'h0616;    16'd11190: out <= 16'h06A4;    16'd11191: out <= 16'h01E6;
    16'd11192: out <= 16'h05EC;    16'd11193: out <= 16'hFF8A;    16'd11194: out <= 16'hFD83;    16'd11195: out <= 16'hFF64;
    16'd11196: out <= 16'h0450;    16'd11197: out <= 16'h02C2;    16'd11198: out <= 16'hFED9;    16'd11199: out <= 16'h0935;
    16'd11200: out <= 16'h054F;    16'd11201: out <= 16'h0387;    16'd11202: out <= 16'h01CF;    16'd11203: out <= 16'h01B2;
    16'd11204: out <= 16'h0250;    16'd11205: out <= 16'h0949;    16'd11206: out <= 16'h066E;    16'd11207: out <= 16'h02B8;
    16'd11208: out <= 16'h0704;    16'd11209: out <= 16'h06E2;    16'd11210: out <= 16'h094F;    16'd11211: out <= 16'h0341;
    16'd11212: out <= 16'h02B9;    16'd11213: out <= 16'h04E8;    16'd11214: out <= 16'h02D8;    16'd11215: out <= 16'h0127;
    16'd11216: out <= 16'h0716;    16'd11217: out <= 16'h0197;    16'd11218: out <= 16'hFF8B;    16'd11219: out <= 16'hFE3F;
    16'd11220: out <= 16'hFF7C;    16'd11221: out <= 16'hFCB9;    16'd11222: out <= 16'h0237;    16'd11223: out <= 16'hF9BF;
    16'd11224: out <= 16'h0187;    16'd11225: out <= 16'hFE72;    16'd11226: out <= 16'hFD94;    16'd11227: out <= 16'hF7C1;
    16'd11228: out <= 16'h02EF;    16'd11229: out <= 16'h04E0;    16'd11230: out <= 16'hFE5E;    16'd11231: out <= 16'hFB19;
    16'd11232: out <= 16'h022B;    16'd11233: out <= 16'hFCD0;    16'd11234: out <= 16'h017A;    16'd11235: out <= 16'h0061;
    16'd11236: out <= 16'hFF48;    16'd11237: out <= 16'h0661;    16'd11238: out <= 16'h0114;    16'd11239: out <= 16'h09DE;
    16'd11240: out <= 16'hF859;    16'd11241: out <= 16'hFBD3;    16'd11242: out <= 16'h03A3;    16'd11243: out <= 16'hFB18;
    16'd11244: out <= 16'hFD31;    16'd11245: out <= 16'hFE98;    16'd11246: out <= 16'hFF37;    16'd11247: out <= 16'h0231;
    16'd11248: out <= 16'hFB38;    16'd11249: out <= 16'hFB12;    16'd11250: out <= 16'hFE8B;    16'd11251: out <= 16'hFF89;
    16'd11252: out <= 16'h004F;    16'd11253: out <= 16'hFEDF;    16'd11254: out <= 16'hFC17;    16'd11255: out <= 16'h02F2;
    16'd11256: out <= 16'h04C7;    16'd11257: out <= 16'h04DD;    16'd11258: out <= 16'hFB16;    16'd11259: out <= 16'h0341;
    16'd11260: out <= 16'h047B;    16'd11261: out <= 16'hF4F3;    16'd11262: out <= 16'hFDCC;    16'd11263: out <= 16'hFBC7;
    16'd11264: out <= 16'h00DB;    16'd11265: out <= 16'h04C7;    16'd11266: out <= 16'h07B6;    16'd11267: out <= 16'hFB8F;
    16'd11268: out <= 16'h03EE;    16'd11269: out <= 16'hFBA5;    16'd11270: out <= 16'h02C3;    16'd11271: out <= 16'h04BD;
    16'd11272: out <= 16'hF592;    16'd11273: out <= 16'hFF02;    16'd11274: out <= 16'h0163;    16'd11275: out <= 16'hFF91;
    16'd11276: out <= 16'hFE18;    16'd11277: out <= 16'hF909;    16'd11278: out <= 16'hFF7C;    16'd11279: out <= 16'hFCE2;
    16'd11280: out <= 16'h0482;    16'd11281: out <= 16'h0012;    16'd11282: out <= 16'hFE2D;    16'd11283: out <= 16'h03F4;
    16'd11284: out <= 16'h0113;    16'd11285: out <= 16'h03DD;    16'd11286: out <= 16'hFDB1;    16'd11287: out <= 16'hFEFC;
    16'd11288: out <= 16'h04E7;    16'd11289: out <= 16'hFA62;    16'd11290: out <= 16'hFC59;    16'd11291: out <= 16'hFF37;
    16'd11292: out <= 16'hFFDC;    16'd11293: out <= 16'hFB15;    16'd11294: out <= 16'hF704;    16'd11295: out <= 16'h013D;
    16'd11296: out <= 16'h00BC;    16'd11297: out <= 16'h0037;    16'd11298: out <= 16'hFEA6;    16'd11299: out <= 16'h054E;
    16'd11300: out <= 16'h0266;    16'd11301: out <= 16'h0028;    16'd11302: out <= 16'h08F9;    16'd11303: out <= 16'h039E;
    16'd11304: out <= 16'h0398;    16'd11305: out <= 16'h023C;    16'd11306: out <= 16'h0222;    16'd11307: out <= 16'h0A60;
    16'd11308: out <= 16'h04C6;    16'd11309: out <= 16'h04AA;    16'd11310: out <= 16'h0827;    16'd11311: out <= 16'h04AD;
    16'd11312: out <= 16'hFC81;    16'd11313: out <= 16'h0454;    16'd11314: out <= 16'h03A5;    16'd11315: out <= 16'h00D8;
    16'd11316: out <= 16'h0318;    16'd11317: out <= 16'h077B;    16'd11318: out <= 16'h06A0;    16'd11319: out <= 16'h00DF;
    16'd11320: out <= 16'h0374;    16'd11321: out <= 16'h018D;    16'd11322: out <= 16'h05F3;    16'd11323: out <= 16'hFF46;
    16'd11324: out <= 16'h0559;    16'd11325: out <= 16'h002A;    16'd11326: out <= 16'h05FC;    16'd11327: out <= 16'h05C5;
    16'd11328: out <= 16'h0848;    16'd11329: out <= 16'h0000;    16'd11330: out <= 16'hFC8D;    16'd11331: out <= 16'h0334;
    16'd11332: out <= 16'h0119;    16'd11333: out <= 16'hFCAA;    16'd11334: out <= 16'h045A;    16'd11335: out <= 16'h0C32;
    16'd11336: out <= 16'h0A04;    16'd11337: out <= 16'hFB97;    16'd11338: out <= 16'h1104;    16'd11339: out <= 16'h0054;
    16'd11340: out <= 16'h0574;    16'd11341: out <= 16'h001F;    16'd11342: out <= 16'h0662;    16'd11343: out <= 16'h0106;
    16'd11344: out <= 16'h0629;    16'd11345: out <= 16'hFE7D;    16'd11346: out <= 16'h0355;    16'd11347: out <= 16'h06FF;
    16'd11348: out <= 16'h03AD;    16'd11349: out <= 16'h0275;    16'd11350: out <= 16'h05A2;    16'd11351: out <= 16'h0797;
    16'd11352: out <= 16'h062D;    16'd11353: out <= 16'h05B9;    16'd11354: out <= 16'h0362;    16'd11355: out <= 16'hFA07;
    16'd11356: out <= 16'h06BF;    16'd11357: out <= 16'h080F;    16'd11358: out <= 16'h03E7;    16'd11359: out <= 16'h08DE;
    16'd11360: out <= 16'h051C;    16'd11361: out <= 16'h067D;    16'd11362: out <= 16'h039E;    16'd11363: out <= 16'hFE2C;
    16'd11364: out <= 16'hFB36;    16'd11365: out <= 16'h037B;    16'd11366: out <= 16'h0550;    16'd11367: out <= 16'hFF3B;
    16'd11368: out <= 16'h0656;    16'd11369: out <= 16'h038F;    16'd11370: out <= 16'h022B;    16'd11371: out <= 16'h022F;
    16'd11372: out <= 16'h0577;    16'd11373: out <= 16'h0749;    16'd11374: out <= 16'hFCF3;    16'd11375: out <= 16'h032F;
    16'd11376: out <= 16'hFC87;    16'd11377: out <= 16'h00D5;    16'd11378: out <= 16'h067C;    16'd11379: out <= 16'h05FC;
    16'd11380: out <= 16'h021F;    16'd11381: out <= 16'h011E;    16'd11382: out <= 16'h032B;    16'd11383: out <= 16'h0082;
    16'd11384: out <= 16'h0465;    16'd11385: out <= 16'h01E0;    16'd11386: out <= 16'hFAD7;    16'd11387: out <= 16'h0455;
    16'd11388: out <= 16'hFE9E;    16'd11389: out <= 16'h03F4;    16'd11390: out <= 16'hFDB5;    16'd11391: out <= 16'hFCD4;
    16'd11392: out <= 16'h0473;    16'd11393: out <= 16'h054A;    16'd11394: out <= 16'h049C;    16'd11395: out <= 16'h0242;
    16'd11396: out <= 16'h054D;    16'd11397: out <= 16'h0326;    16'd11398: out <= 16'hFFAD;    16'd11399: out <= 16'h0009;
    16'd11400: out <= 16'h0529;    16'd11401: out <= 16'hFF62;    16'd11402: out <= 16'h0261;    16'd11403: out <= 16'h0800;
    16'd11404: out <= 16'h02D9;    16'd11405: out <= 16'h0726;    16'd11406: out <= 16'h0106;    16'd11407: out <= 16'h0257;
    16'd11408: out <= 16'h0830;    16'd11409: out <= 16'h01D7;    16'd11410: out <= 16'h028E;    16'd11411: out <= 16'hFE27;
    16'd11412: out <= 16'h017B;    16'd11413: out <= 16'h084D;    16'd11414: out <= 16'h01F3;    16'd11415: out <= 16'h0252;
    16'd11416: out <= 16'h0839;    16'd11417: out <= 16'h0735;    16'd11418: out <= 16'hFE0B;    16'd11419: out <= 16'h0698;
    16'd11420: out <= 16'h00C8;    16'd11421: out <= 16'h0288;    16'd11422: out <= 16'h0310;    16'd11423: out <= 16'h0144;
    16'd11424: out <= 16'h0107;    16'd11425: out <= 16'h04C9;    16'd11426: out <= 16'h0201;    16'd11427: out <= 16'h055B;
    16'd11428: out <= 16'hFF48;    16'd11429: out <= 16'h048A;    16'd11430: out <= 16'h06EA;    16'd11431: out <= 16'h0545;
    16'd11432: out <= 16'h0585;    16'd11433: out <= 16'h047B;    16'd11434: out <= 16'h06C9;    16'd11435: out <= 16'h0916;
    16'd11436: out <= 16'h0610;    16'd11437: out <= 16'h0873;    16'd11438: out <= 16'h0E95;    16'd11439: out <= 16'h0193;
    16'd11440: out <= 16'h03D4;    16'd11441: out <= 16'hFE7E;    16'd11442: out <= 16'h020E;    16'd11443: out <= 16'h0354;
    16'd11444: out <= 16'h0774;    16'd11445: out <= 16'h01C9;    16'd11446: out <= 16'h09B9;    16'd11447: out <= 16'hFF91;
    16'd11448: out <= 16'h050C;    16'd11449: out <= 16'h032B;    16'd11450: out <= 16'h0451;    16'd11451: out <= 16'hFDA2;
    16'd11452: out <= 16'h0C97;    16'd11453: out <= 16'h09C9;    16'd11454: out <= 16'h03F4;    16'd11455: out <= 16'hFF58;
    16'd11456: out <= 16'h061B;    16'd11457: out <= 16'h04EA;    16'd11458: out <= 16'h04D9;    16'd11459: out <= 16'h0493;
    16'd11460: out <= 16'h07CA;    16'd11461: out <= 16'h03DE;    16'd11462: out <= 16'h0882;    16'd11463: out <= 16'h0DD6;
    16'd11464: out <= 16'h0650;    16'd11465: out <= 16'h074A;    16'd11466: out <= 16'h03B7;    16'd11467: out <= 16'h0955;
    16'd11468: out <= 16'h0151;    16'd11469: out <= 16'h0C69;    16'd11470: out <= 16'h0499;    16'd11471: out <= 16'h06C6;
    16'd11472: out <= 16'h02D8;    16'd11473: out <= 16'h0565;    16'd11474: out <= 16'h0248;    16'd11475: out <= 16'h0379;
    16'd11476: out <= 16'h04D6;    16'd11477: out <= 16'hFA69;    16'd11478: out <= 16'h023C;    16'd11479: out <= 16'h0752;
    16'd11480: out <= 16'hFAAD;    16'd11481: out <= 16'h06E5;    16'd11482: out <= 16'h03BD;    16'd11483: out <= 16'h0314;
    16'd11484: out <= 16'h02C5;    16'd11485: out <= 16'h0392;    16'd11486: out <= 16'hFA2C;    16'd11487: out <= 16'h0092;
    16'd11488: out <= 16'h0646;    16'd11489: out <= 16'h03D0;    16'd11490: out <= 16'hFC18;    16'd11491: out <= 16'hFAD7;
    16'd11492: out <= 16'hFA50;    16'd11493: out <= 16'h03BF;    16'd11494: out <= 16'hFD6A;    16'd11495: out <= 16'h04C5;
    16'd11496: out <= 16'hFCD0;    16'd11497: out <= 16'hFF3B;    16'd11498: out <= 16'hFED8;    16'd11499: out <= 16'hFFE7;
    16'd11500: out <= 16'h0479;    16'd11501: out <= 16'hF97F;    16'd11502: out <= 16'hFFD1;    16'd11503: out <= 16'h03F2;
    16'd11504: out <= 16'hFE30;    16'd11505: out <= 16'h0003;    16'd11506: out <= 16'h0248;    16'd11507: out <= 16'h0688;
    16'd11508: out <= 16'hFB9F;    16'd11509: out <= 16'h007D;    16'd11510: out <= 16'hF881;    16'd11511: out <= 16'hFAF8;
    16'd11512: out <= 16'hFD0D;    16'd11513: out <= 16'h0556;    16'd11514: out <= 16'h0224;    16'd11515: out <= 16'h076B;
    16'd11516: out <= 16'hFCC5;    16'd11517: out <= 16'h01A3;    16'd11518: out <= 16'h0485;    16'd11519: out <= 16'hFF44;
    16'd11520: out <= 16'h07CA;    16'd11521: out <= 16'h0802;    16'd11522: out <= 16'hFC66;    16'd11523: out <= 16'h0176;
    16'd11524: out <= 16'h01BB;    16'd11525: out <= 16'h044B;    16'd11526: out <= 16'hFD91;    16'd11527: out <= 16'hFCFD;
    16'd11528: out <= 16'h08BA;    16'd11529: out <= 16'h0024;    16'd11530: out <= 16'hF6C3;    16'd11531: out <= 16'hFEF8;
    16'd11532: out <= 16'h05E4;    16'd11533: out <= 16'h00C3;    16'd11534: out <= 16'hFDB2;    16'd11535: out <= 16'h036F;
    16'd11536: out <= 16'hFB07;    16'd11537: out <= 16'hF8C5;    16'd11538: out <= 16'h028C;    16'd11539: out <= 16'hF6D5;
    16'd11540: out <= 16'h009D;    16'd11541: out <= 16'hFD7C;    16'd11542: out <= 16'h010B;    16'd11543: out <= 16'h021A;
    16'd11544: out <= 16'hF908;    16'd11545: out <= 16'hFD3D;    16'd11546: out <= 16'h0525;    16'd11547: out <= 16'hFC29;
    16'd11548: out <= 16'hFEB6;    16'd11549: out <= 16'hFF30;    16'd11550: out <= 16'h0441;    16'd11551: out <= 16'h0114;
    16'd11552: out <= 16'hFE42;    16'd11553: out <= 16'h02C1;    16'd11554: out <= 16'h0040;    16'd11555: out <= 16'h027E;
    16'd11556: out <= 16'h010C;    16'd11557: out <= 16'h053C;    16'd11558: out <= 16'h04AC;    16'd11559: out <= 16'h0189;
    16'd11560: out <= 16'hFD5D;    16'd11561: out <= 16'h0039;    16'd11562: out <= 16'h07E9;    16'd11563: out <= 16'h0362;
    16'd11564: out <= 16'hFE4E;    16'd11565: out <= 16'h06C1;    16'd11566: out <= 16'h074F;    16'd11567: out <= 16'hFD48;
    16'd11568: out <= 16'hFFD2;    16'd11569: out <= 16'h031C;    16'd11570: out <= 16'h0223;    16'd11571: out <= 16'h0883;
    16'd11572: out <= 16'h055C;    16'd11573: out <= 16'h0D27;    16'd11574: out <= 16'h05D7;    16'd11575: out <= 16'h074F;
    16'd11576: out <= 16'h0190;    16'd11577: out <= 16'h0743;    16'd11578: out <= 16'h04AA;    16'd11579: out <= 16'hFF89;
    16'd11580: out <= 16'hFF94;    16'd11581: out <= 16'h07C6;    16'd11582: out <= 16'h05AF;    16'd11583: out <= 16'h07EB;
    16'd11584: out <= 16'h026C;    16'd11585: out <= 16'h02AC;    16'd11586: out <= 16'h064B;    16'd11587: out <= 16'h07A5;
    16'd11588: out <= 16'h02FC;    16'd11589: out <= 16'hFCE8;    16'd11590: out <= 16'h0006;    16'd11591: out <= 16'h09EA;
    16'd11592: out <= 16'h041D;    16'd11593: out <= 16'h039E;    16'd11594: out <= 16'h0736;    16'd11595: out <= 16'hFEF6;
    16'd11596: out <= 16'h0229;    16'd11597: out <= 16'h008C;    16'd11598: out <= 16'h03AD;    16'd11599: out <= 16'h0902;
    16'd11600: out <= 16'h0003;    16'd11601: out <= 16'h00CE;    16'd11602: out <= 16'h03DF;    16'd11603: out <= 16'hFF31;
    16'd11604: out <= 16'h0630;    16'd11605: out <= 16'h0BB0;    16'd11606: out <= 16'h0CEC;    16'd11607: out <= 16'h0441;
    16'd11608: out <= 16'h09EB;    16'd11609: out <= 16'h02BC;    16'd11610: out <= 16'h020C;    16'd11611: out <= 16'h019E;
    16'd11612: out <= 16'hFD49;    16'd11613: out <= 16'h06CA;    16'd11614: out <= 16'h03C1;    16'd11615: out <= 16'hFE27;
    16'd11616: out <= 16'h0335;    16'd11617: out <= 16'h08A5;    16'd11618: out <= 16'h08B5;    16'd11619: out <= 16'h040B;
    16'd11620: out <= 16'h0D5A;    16'd11621: out <= 16'h01F0;    16'd11622: out <= 16'h0437;    16'd11623: out <= 16'hFCAE;
    16'd11624: out <= 16'h0511;    16'd11625: out <= 16'h0812;    16'd11626: out <= 16'h0843;    16'd11627: out <= 16'h05D5;
    16'd11628: out <= 16'h009C;    16'd11629: out <= 16'h0E4F;    16'd11630: out <= 16'h0C99;    16'd11631: out <= 16'h005A;
    16'd11632: out <= 16'h0198;    16'd11633: out <= 16'h0021;    16'd11634: out <= 16'h064F;    16'd11635: out <= 16'hFF29;
    16'd11636: out <= 16'h02D2;    16'd11637: out <= 16'h080F;    16'd11638: out <= 16'h06D6;    16'd11639: out <= 16'hFDD8;
    16'd11640: out <= 16'h00FF;    16'd11641: out <= 16'h063B;    16'd11642: out <= 16'h0031;    16'd11643: out <= 16'h0457;
    16'd11644: out <= 16'h07AF;    16'd11645: out <= 16'h07DD;    16'd11646: out <= 16'h0A58;    16'd11647: out <= 16'h0105;
    16'd11648: out <= 16'h04B5;    16'd11649: out <= 16'h0309;    16'd11650: out <= 16'h0C03;    16'd11651: out <= 16'h0615;
    16'd11652: out <= 16'h08D3;    16'd11653: out <= 16'hFF16;    16'd11654: out <= 16'hFDF9;    16'd11655: out <= 16'hFFB5;
    16'd11656: out <= 16'hFD03;    16'd11657: out <= 16'h0621;    16'd11658: out <= 16'h0694;    16'd11659: out <= 16'h0391;
    16'd11660: out <= 16'h007A;    16'd11661: out <= 16'h048F;    16'd11662: out <= 16'hFD70;    16'd11663: out <= 16'h016C;
    16'd11664: out <= 16'h070B;    16'd11665: out <= 16'h011C;    16'd11666: out <= 16'h0372;    16'd11667: out <= 16'h06D9;
    16'd11668: out <= 16'h0C23;    16'd11669: out <= 16'h0422;    16'd11670: out <= 16'h003B;    16'd11671: out <= 16'h0583;
    16'd11672: out <= 16'h04EB;    16'd11673: out <= 16'h07F9;    16'd11674: out <= 16'h025E;    16'd11675: out <= 16'h0310;
    16'd11676: out <= 16'hFCF2;    16'd11677: out <= 16'hFF76;    16'd11678: out <= 16'h02E7;    16'd11679: out <= 16'h021E;
    16'd11680: out <= 16'h0173;    16'd11681: out <= 16'h0753;    16'd11682: out <= 16'h0796;    16'd11683: out <= 16'h04E2;
    16'd11684: out <= 16'h006B;    16'd11685: out <= 16'hFE52;    16'd11686: out <= 16'hFDD9;    16'd11687: out <= 16'h04DE;
    16'd11688: out <= 16'h0889;    16'd11689: out <= 16'h054F;    16'd11690: out <= 16'h0698;    16'd11691: out <= 16'h007A;
    16'd11692: out <= 16'h0163;    16'd11693: out <= 16'hFE26;    16'd11694: out <= 16'hFB79;    16'd11695: out <= 16'hF92C;
    16'd11696: out <= 16'hFFA7;    16'd11697: out <= 16'h06E6;    16'd11698: out <= 16'h0065;    16'd11699: out <= 16'h03D8;
    16'd11700: out <= 16'h02B8;    16'd11701: out <= 16'h0821;    16'd11702: out <= 16'h09AE;    16'd11703: out <= 16'h0346;
    16'd11704: out <= 16'h030D;    16'd11705: out <= 16'h06D6;    16'd11706: out <= 16'h0626;    16'd11707: out <= 16'h0640;
    16'd11708: out <= 16'hF9D3;    16'd11709: out <= 16'h00A9;    16'd11710: out <= 16'h032E;    16'd11711: out <= 16'h069A;
    16'd11712: out <= 16'h05C5;    16'd11713: out <= 16'h03C0;    16'd11714: out <= 16'hFF77;    16'd11715: out <= 16'h07E4;
    16'd11716: out <= 16'h0091;    16'd11717: out <= 16'hFD10;    16'd11718: out <= 16'h0C35;    16'd11719: out <= 16'h02CF;
    16'd11720: out <= 16'h044D;    16'd11721: out <= 16'hFEBE;    16'd11722: out <= 16'h06BF;    16'd11723: out <= 16'h0964;
    16'd11724: out <= 16'h0A31;    16'd11725: out <= 16'h02DD;    16'd11726: out <= 16'h01B5;    16'd11727: out <= 16'h04AB;
    16'd11728: out <= 16'h017E;    16'd11729: out <= 16'h02D5;    16'd11730: out <= 16'h09D7;    16'd11731: out <= 16'h051E;
    16'd11732: out <= 16'h013D;    16'd11733: out <= 16'hFF21;    16'd11734: out <= 16'h00AD;    16'd11735: out <= 16'h03A5;
    16'd11736: out <= 16'h0044;    16'd11737: out <= 16'h02BE;    16'd11738: out <= 16'hFD3E;    16'd11739: out <= 16'h03B7;
    16'd11740: out <= 16'hFE59;    16'd11741: out <= 16'h01F6;    16'd11742: out <= 16'h0146;    16'd11743: out <= 16'hFA7B;
    16'd11744: out <= 16'hFD5B;    16'd11745: out <= 16'h0382;    16'd11746: out <= 16'h02B9;    16'd11747: out <= 16'h00CE;
    16'd11748: out <= 16'hF864;    16'd11749: out <= 16'hFF9F;    16'd11750: out <= 16'h01BC;    16'd11751: out <= 16'h03A2;
    16'd11752: out <= 16'hFDB8;    16'd11753: out <= 16'hFA00;    16'd11754: out <= 16'hFF67;    16'd11755: out <= 16'hFEB8;
    16'd11756: out <= 16'hFF2A;    16'd11757: out <= 16'h04EF;    16'd11758: out <= 16'h033F;    16'd11759: out <= 16'h0005;
    16'd11760: out <= 16'hFDB3;    16'd11761: out <= 16'h00FB;    16'd11762: out <= 16'hFE9C;    16'd11763: out <= 16'hFE49;
    16'd11764: out <= 16'hFE81;    16'd11765: out <= 16'h00C9;    16'd11766: out <= 16'h03F5;    16'd11767: out <= 16'hFF99;
    16'd11768: out <= 16'h00C3;    16'd11769: out <= 16'h05B6;    16'd11770: out <= 16'hFC29;    16'd11771: out <= 16'hFCC4;
    16'd11772: out <= 16'hFCFF;    16'd11773: out <= 16'h04DB;    16'd11774: out <= 16'hFEA0;    16'd11775: out <= 16'h06BC;
    16'd11776: out <= 16'hFDCB;    16'd11777: out <= 16'hFE65;    16'd11778: out <= 16'h04F9;    16'd11779: out <= 16'h0015;
    16'd11780: out <= 16'h04C1;    16'd11781: out <= 16'h079B;    16'd11782: out <= 16'hFEBB;    16'd11783: out <= 16'hFEBA;
    16'd11784: out <= 16'hFFED;    16'd11785: out <= 16'hFC4A;    16'd11786: out <= 16'hFB62;    16'd11787: out <= 16'hF64B;
    16'd11788: out <= 16'h007B;    16'd11789: out <= 16'h0013;    16'd11790: out <= 16'h0395;    16'd11791: out <= 16'hFC5F;
    16'd11792: out <= 16'h028C;    16'd11793: out <= 16'hFF3A;    16'd11794: out <= 16'h0392;    16'd11795: out <= 16'hFEFE;
    16'd11796: out <= 16'h0780;    16'd11797: out <= 16'hFBF1;    16'd11798: out <= 16'h03B5;    16'd11799: out <= 16'hF820;
    16'd11800: out <= 16'h018D;    16'd11801: out <= 16'hF713;    16'd11802: out <= 16'hFFF2;    16'd11803: out <= 16'h02F7;
    16'd11804: out <= 16'h027E;    16'd11805: out <= 16'hFF22;    16'd11806: out <= 16'h00E6;    16'd11807: out <= 16'hFF30;
    16'd11808: out <= 16'hFEC3;    16'd11809: out <= 16'hFD95;    16'd11810: out <= 16'h0419;    16'd11811: out <= 16'h0225;
    16'd11812: out <= 16'h0492;    16'd11813: out <= 16'h0595;    16'd11814: out <= 16'h0170;    16'd11815: out <= 16'h01BA;
    16'd11816: out <= 16'h0A6F;    16'd11817: out <= 16'h0BA4;    16'd11818: out <= 16'h0290;    16'd11819: out <= 16'h0D5E;
    16'd11820: out <= 16'hFF14;    16'd11821: out <= 16'h0690;    16'd11822: out <= 16'hFBE6;    16'd11823: out <= 16'hFD79;
    16'd11824: out <= 16'h03B3;    16'd11825: out <= 16'h01CE;    16'd11826: out <= 16'h0237;    16'd11827: out <= 16'h0833;
    16'd11828: out <= 16'h0592;    16'd11829: out <= 16'h01C2;    16'd11830: out <= 16'hFDF9;    16'd11831: out <= 16'h0B00;
    16'd11832: out <= 16'hFD0E;    16'd11833: out <= 16'h011F;    16'd11834: out <= 16'h02A5;    16'd11835: out <= 16'h03AC;
    16'd11836: out <= 16'h09A1;    16'd11837: out <= 16'h005A;    16'd11838: out <= 16'h0587;    16'd11839: out <= 16'hFE67;
    16'd11840: out <= 16'h075A;    16'd11841: out <= 16'h0384;    16'd11842: out <= 16'hFD39;    16'd11843: out <= 16'h1138;
    16'd11844: out <= 16'h091B;    16'd11845: out <= 16'hFA26;    16'd11846: out <= 16'h002A;    16'd11847: out <= 16'h0202;
    16'd11848: out <= 16'h024F;    16'd11849: out <= 16'h00A6;    16'd11850: out <= 16'h07CB;    16'd11851: out <= 16'h0CFF;
    16'd11852: out <= 16'h0485;    16'd11853: out <= 16'h070E;    16'd11854: out <= 16'h0088;    16'd11855: out <= 16'h04D8;
    16'd11856: out <= 16'h0154;    16'd11857: out <= 16'h0933;    16'd11858: out <= 16'h0682;    16'd11859: out <= 16'h02C3;
    16'd11860: out <= 16'h0AFF;    16'd11861: out <= 16'h0699;    16'd11862: out <= 16'h01D7;    16'd11863: out <= 16'h026C;
    16'd11864: out <= 16'h0326;    16'd11865: out <= 16'h03E8;    16'd11866: out <= 16'h041C;    16'd11867: out <= 16'h00BE;
    16'd11868: out <= 16'h0275;    16'd11869: out <= 16'h01E2;    16'd11870: out <= 16'h05BE;    16'd11871: out <= 16'hFF4E;
    16'd11872: out <= 16'h00BA;    16'd11873: out <= 16'h047B;    16'd11874: out <= 16'h0852;    16'd11875: out <= 16'h0062;
    16'd11876: out <= 16'h0680;    16'd11877: out <= 16'h0E4F;    16'd11878: out <= 16'h00C4;    16'd11879: out <= 16'h001F;
    16'd11880: out <= 16'h07C8;    16'd11881: out <= 16'h081B;    16'd11882: out <= 16'h0AE4;    16'd11883: out <= 16'h0100;
    16'd11884: out <= 16'h0743;    16'd11885: out <= 16'h00CA;    16'd11886: out <= 16'hFCB5;    16'd11887: out <= 16'h0750;
    16'd11888: out <= 16'h0029;    16'd11889: out <= 16'h0476;    16'd11890: out <= 16'h0334;    16'd11891: out <= 16'h0557;
    16'd11892: out <= 16'h02AB;    16'd11893: out <= 16'h083F;    16'd11894: out <= 16'h06FE;    16'd11895: out <= 16'h04D3;
    16'd11896: out <= 16'hFFB5;    16'd11897: out <= 16'h09A5;    16'd11898: out <= 16'h0D5D;    16'd11899: out <= 16'h024A;
    16'd11900: out <= 16'h0235;    16'd11901: out <= 16'hFA97;    16'd11902: out <= 16'h05FC;    16'd11903: out <= 16'h0589;
    16'd11904: out <= 16'h0239;    16'd11905: out <= 16'h016A;    16'd11906: out <= 16'h0895;    16'd11907: out <= 16'hFD17;
    16'd11908: out <= 16'hFFB1;    16'd11909: out <= 16'hFD5C;    16'd11910: out <= 16'h0141;    16'd11911: out <= 16'h0C8C;
    16'd11912: out <= 16'hFCD0;    16'd11913: out <= 16'h0492;    16'd11914: out <= 16'hF7C8;    16'd11915: out <= 16'h039C;
    16'd11916: out <= 16'h00C8;    16'd11917: out <= 16'h0424;    16'd11918: out <= 16'h0C08;    16'd11919: out <= 16'h02DB;
    16'd11920: out <= 16'h0A54;    16'd11921: out <= 16'h0A4A;    16'd11922: out <= 16'h01CC;    16'd11923: out <= 16'h08D2;
    16'd11924: out <= 16'h037C;    16'd11925: out <= 16'h056D;    16'd11926: out <= 16'hFE10;    16'd11927: out <= 16'h08D4;
    16'd11928: out <= 16'h09BC;    16'd11929: out <= 16'h0124;    16'd11930: out <= 16'h0362;    16'd11931: out <= 16'h04C8;
    16'd11932: out <= 16'hFAF4;    16'd11933: out <= 16'h0497;    16'd11934: out <= 16'h0441;    16'd11935: out <= 16'h0984;
    16'd11936: out <= 16'h09E6;    16'd11937: out <= 16'h05F8;    16'd11938: out <= 16'h02F1;    16'd11939: out <= 16'hFEE7;
    16'd11940: out <= 16'hFFEC;    16'd11941: out <= 16'h01D2;    16'd11942: out <= 16'h0255;    16'd11943: out <= 16'h06C8;
    16'd11944: out <= 16'h01E4;    16'd11945: out <= 16'h02BC;    16'd11946: out <= 16'h03AC;    16'd11947: out <= 16'hFE34;
    16'd11948: out <= 16'hFC9B;    16'd11949: out <= 16'h0488;    16'd11950: out <= 16'h03B0;    16'd11951: out <= 16'h0338;
    16'd11952: out <= 16'h06FC;    16'd11953: out <= 16'h0A28;    16'd11954: out <= 16'h0187;    16'd11955: out <= 16'h021C;
    16'd11956: out <= 16'h0617;    16'd11957: out <= 16'h06B0;    16'd11958: out <= 16'hFE29;    16'd11959: out <= 16'hFDA5;
    16'd11960: out <= 16'h0557;    16'd11961: out <= 16'h0808;    16'd11962: out <= 16'hFE95;    16'd11963: out <= 16'h031C;
    16'd11964: out <= 16'h04AA;    16'd11965: out <= 16'h040B;    16'd11966: out <= 16'h0276;    16'd11967: out <= 16'h024D;
    16'd11968: out <= 16'h0E4E;    16'd11969: out <= 16'h04E8;    16'd11970: out <= 16'h022F;    16'd11971: out <= 16'h0374;
    16'd11972: out <= 16'hFF96;    16'd11973: out <= 16'h02E4;    16'd11974: out <= 16'h00E0;    16'd11975: out <= 16'h0698;
    16'd11976: out <= 16'h0A2F;    16'd11977: out <= 16'hFF94;    16'd11978: out <= 16'h07FF;    16'd11979: out <= 16'h0568;
    16'd11980: out <= 16'h050F;    16'd11981: out <= 16'h0613;    16'd11982: out <= 16'h02BE;    16'd11983: out <= 16'h0150;
    16'd11984: out <= 16'h0304;    16'd11985: out <= 16'h09F5;    16'd11986: out <= 16'h057D;    16'd11987: out <= 16'h0497;
    16'd11988: out <= 16'h00AE;    16'd11989: out <= 16'hF8FE;    16'd11990: out <= 16'hFAE1;    16'd11991: out <= 16'hFC1A;
    16'd11992: out <= 16'hFBFF;    16'd11993: out <= 16'hFDBF;    16'd11994: out <= 16'hFC40;    16'd11995: out <= 16'h0386;
    16'd11996: out <= 16'hFEF8;    16'd11997: out <= 16'h045F;    16'd11998: out <= 16'h0308;    16'd11999: out <= 16'hFD43;
    16'd12000: out <= 16'h0357;    16'd12001: out <= 16'h04B4;    16'd12002: out <= 16'hFED9;    16'd12003: out <= 16'hFCE3;
    16'd12004: out <= 16'h0095;    16'd12005: out <= 16'h05DB;    16'd12006: out <= 16'hF963;    16'd12007: out <= 16'h02D9;
    16'd12008: out <= 16'hFF44;    16'd12009: out <= 16'h0447;    16'd12010: out <= 16'hFF8C;    16'd12011: out <= 16'hFCC6;
    16'd12012: out <= 16'h0062;    16'd12013: out <= 16'h0190;    16'd12014: out <= 16'h037E;    16'd12015: out <= 16'h05A6;
    16'd12016: out <= 16'hFFA4;    16'd12017: out <= 16'h0464;    16'd12018: out <= 16'hFF2B;    16'd12019: out <= 16'h00C9;
    16'd12020: out <= 16'h0188;    16'd12021: out <= 16'h08FF;    16'd12022: out <= 16'hFEFB;    16'd12023: out <= 16'hFF62;
    16'd12024: out <= 16'hFF1A;    16'd12025: out <= 16'h009F;    16'd12026: out <= 16'h0161;    16'd12027: out <= 16'hFC3D;
    16'd12028: out <= 16'hFC9B;    16'd12029: out <= 16'h010B;    16'd12030: out <= 16'hFDF1;    16'd12031: out <= 16'h0178;
    16'd12032: out <= 16'hFABD;    16'd12033: out <= 16'hF6A0;    16'd12034: out <= 16'h068C;    16'd12035: out <= 16'hFF86;
    16'd12036: out <= 16'hFFD1;    16'd12037: out <= 16'hF807;    16'd12038: out <= 16'h01C0;    16'd12039: out <= 16'h03AC;
    16'd12040: out <= 16'h032F;    16'd12041: out <= 16'hFD73;    16'd12042: out <= 16'h018C;    16'd12043: out <= 16'hFDAF;
    16'd12044: out <= 16'hFC74;    16'd12045: out <= 16'h01AA;    16'd12046: out <= 16'h02D7;    16'd12047: out <= 16'h014B;
    16'd12048: out <= 16'h01F8;    16'd12049: out <= 16'hFEA4;    16'd12050: out <= 16'hFCEB;    16'd12051: out <= 16'h02AA;
    16'd12052: out <= 16'hFD2C;    16'd12053: out <= 16'hFAF0;    16'd12054: out <= 16'hFE33;    16'd12055: out <= 16'hF8E2;
    16'd12056: out <= 16'h0833;    16'd12057: out <= 16'h05F6;    16'd12058: out <= 16'hFFFB;    16'd12059: out <= 16'h0151;
    16'd12060: out <= 16'h0092;    16'd12061: out <= 16'h0132;    16'd12062: out <= 16'hFE25;    16'd12063: out <= 16'h03FB;
    16'd12064: out <= 16'h04C8;    16'd12065: out <= 16'hFFBE;    16'd12066: out <= 16'hFD8D;    16'd12067: out <= 16'h03AE;
    16'd12068: out <= 16'hFE73;    16'd12069: out <= 16'hFF2B;    16'd12070: out <= 16'h0606;    16'd12071: out <= 16'h0844;
    16'd12072: out <= 16'hFEFF;    16'd12073: out <= 16'h0870;    16'd12074: out <= 16'h0B6A;    16'd12075: out <= 16'h023A;
    16'd12076: out <= 16'h0721;    16'd12077: out <= 16'h0460;    16'd12078: out <= 16'h05E7;    16'd12079: out <= 16'h060A;
    16'd12080: out <= 16'hF5C2;    16'd12081: out <= 16'h036D;    16'd12082: out <= 16'h0066;    16'd12083: out <= 16'hFE48;
    16'd12084: out <= 16'h05B8;    16'd12085: out <= 16'h0BAF;    16'd12086: out <= 16'h09A6;    16'd12087: out <= 16'h055A;
    16'd12088: out <= 16'h0418;    16'd12089: out <= 16'h0243;    16'd12090: out <= 16'h00D9;    16'd12091: out <= 16'h0882;
    16'd12092: out <= 16'h08C8;    16'd12093: out <= 16'h004E;    16'd12094: out <= 16'h086F;    16'd12095: out <= 16'h01F5;
    16'd12096: out <= 16'h02DE;    16'd12097: out <= 16'h04F7;    16'd12098: out <= 16'h038E;    16'd12099: out <= 16'h073C;
    16'd12100: out <= 16'h0343;    16'd12101: out <= 16'h093F;    16'd12102: out <= 16'h00CE;    16'd12103: out <= 16'hFDF0;
    16'd12104: out <= 16'h0304;    16'd12105: out <= 16'h0539;    16'd12106: out <= 16'h05D9;    16'd12107: out <= 16'hFFA4;
    16'd12108: out <= 16'h0A92;    16'd12109: out <= 16'h0213;    16'd12110: out <= 16'h0618;    16'd12111: out <= 16'h0104;
    16'd12112: out <= 16'h02DC;    16'd12113: out <= 16'h053D;    16'd12114: out <= 16'hFA91;    16'd12115: out <= 16'h0855;
    16'd12116: out <= 16'h046E;    16'd12117: out <= 16'h0472;    16'd12118: out <= 16'h0453;    16'd12119: out <= 16'h03A9;
    16'd12120: out <= 16'h0857;    16'd12121: out <= 16'h0514;    16'd12122: out <= 16'h092E;    16'd12123: out <= 16'h06DE;
    16'd12124: out <= 16'h0018;    16'd12125: out <= 16'h03A7;    16'd12126: out <= 16'hFE2C;    16'd12127: out <= 16'h03F9;
    16'd12128: out <= 16'hFEF5;    16'd12129: out <= 16'h04F7;    16'd12130: out <= 16'h07B7;    16'd12131: out <= 16'h04C4;
    16'd12132: out <= 16'h0303;    16'd12133: out <= 16'h088B;    16'd12134: out <= 16'h07AE;    16'd12135: out <= 16'h03E7;
    16'd12136: out <= 16'h0683;    16'd12137: out <= 16'h070F;    16'd12138: out <= 16'h0258;    16'd12139: out <= 16'h041B;
    16'd12140: out <= 16'hFF52;    16'd12141: out <= 16'h06E1;    16'd12142: out <= 16'h0A9D;    16'd12143: out <= 16'h0015;
    16'd12144: out <= 16'h012D;    16'd12145: out <= 16'h09F4;    16'd12146: out <= 16'h04F6;    16'd12147: out <= 16'h0945;
    16'd12148: out <= 16'hFB93;    16'd12149: out <= 16'hFC42;    16'd12150: out <= 16'h0A79;    16'd12151: out <= 16'h003F;
    16'd12152: out <= 16'h0106;    16'd12153: out <= 16'h01AC;    16'd12154: out <= 16'h074D;    16'd12155: out <= 16'h0374;
    16'd12156: out <= 16'h0B47;    16'd12157: out <= 16'h0897;    16'd12158: out <= 16'h09A8;    16'd12159: out <= 16'h08E5;
    16'd12160: out <= 16'hFD3C;    16'd12161: out <= 16'h052B;    16'd12162: out <= 16'h0653;    16'd12163: out <= 16'h02CE;
    16'd12164: out <= 16'h02BC;    16'd12165: out <= 16'h0020;    16'd12166: out <= 16'h00FC;    16'd12167: out <= 16'h05F8;
    16'd12168: out <= 16'h016C;    16'd12169: out <= 16'h0391;    16'd12170: out <= 16'h00F1;    16'd12171: out <= 16'h0316;
    16'd12172: out <= 16'hFDA0;    16'd12173: out <= 16'h0085;    16'd12174: out <= 16'hFF2D;    16'd12175: out <= 16'h023A;
    16'd12176: out <= 16'h0A50;    16'd12177: out <= 16'hFBA3;    16'd12178: out <= 16'h00AE;    16'd12179: out <= 16'h002C;
    16'd12180: out <= 16'h04C7;    16'd12181: out <= 16'h0671;    16'd12182: out <= 16'h093B;    16'd12183: out <= 16'h08A2;
    16'd12184: out <= 16'hFFA4;    16'd12185: out <= 16'h0189;    16'd12186: out <= 16'hFC19;    16'd12187: out <= 16'h04A4;
    16'd12188: out <= 16'h01EA;    16'd12189: out <= 16'hFF8D;    16'd12190: out <= 16'h0547;    16'd12191: out <= 16'h0386;
    16'd12192: out <= 16'h00C3;    16'd12193: out <= 16'h01F1;    16'd12194: out <= 16'h0430;    16'd12195: out <= 16'hFBDA;
    16'd12196: out <= 16'h07B4;    16'd12197: out <= 16'hFE3C;    16'd12198: out <= 16'h068D;    16'd12199: out <= 16'h0004;
    16'd12200: out <= 16'h0200;    16'd12201: out <= 16'h051D;    16'd12202: out <= 16'h0918;    16'd12203: out <= 16'h083E;
    16'd12204: out <= 16'h06DB;    16'd12205: out <= 16'hFFEF;    16'd12206: out <= 16'h0871;    16'd12207: out <= 16'h0773;
    16'd12208: out <= 16'hFFE7;    16'd12209: out <= 16'h05D3;    16'd12210: out <= 16'h0035;    16'd12211: out <= 16'h01E9;
    16'd12212: out <= 16'h00C4;    16'd12213: out <= 16'h0550;    16'd12214: out <= 16'h0356;    16'd12215: out <= 16'h03A0;
    16'd12216: out <= 16'h0491;    16'd12217: out <= 16'h0581;    16'd12218: out <= 16'h0277;    16'd12219: out <= 16'h01A4;
    16'd12220: out <= 16'h0082;    16'd12221: out <= 16'hFFD7;    16'd12222: out <= 16'h045A;    16'd12223: out <= 16'h0673;
    16'd12224: out <= 16'h0325;    16'd12225: out <= 16'h04D3;    16'd12226: out <= 16'h05C8;    16'd12227: out <= 16'h0567;
    16'd12228: out <= 16'h00FC;    16'd12229: out <= 16'h036B;    16'd12230: out <= 16'hFF2F;    16'd12231: out <= 16'hFFBA;
    16'd12232: out <= 16'h024F;    16'd12233: out <= 16'h03A8;    16'd12234: out <= 16'h0463;    16'd12235: out <= 16'h05FD;
    16'd12236: out <= 16'h04F1;    16'd12237: out <= 16'h0329;    16'd12238: out <= 16'h0817;    16'd12239: out <= 16'h0345;
    16'd12240: out <= 16'h09C1;    16'd12241: out <= 16'h03FE;    16'd12242: out <= 16'hFE9C;    16'd12243: out <= 16'h0325;
    16'd12244: out <= 16'h0462;    16'd12245: out <= 16'h059D;    16'd12246: out <= 16'hFE38;    16'd12247: out <= 16'hFBC5;
    16'd12248: out <= 16'hFB74;    16'd12249: out <= 16'hFF4B;    16'd12250: out <= 16'h0805;    16'd12251: out <= 16'h0396;
    16'd12252: out <= 16'hFECF;    16'd12253: out <= 16'hFF22;    16'd12254: out <= 16'hFBA9;    16'd12255: out <= 16'hFD64;
    16'd12256: out <= 16'h021E;    16'd12257: out <= 16'hF84E;    16'd12258: out <= 16'h0313;    16'd12259: out <= 16'h0773;
    16'd12260: out <= 16'h01FC;    16'd12261: out <= 16'h0510;    16'd12262: out <= 16'h00BC;    16'd12263: out <= 16'hFAEE;
    16'd12264: out <= 16'h0159;    16'd12265: out <= 16'hFE8C;    16'd12266: out <= 16'hFFFD;    16'd12267: out <= 16'h0136;
    16'd12268: out <= 16'h06CD;    16'd12269: out <= 16'h0301;    16'd12270: out <= 16'h00CE;    16'd12271: out <= 16'h0332;
    16'd12272: out <= 16'h083D;    16'd12273: out <= 16'hFD7B;    16'd12274: out <= 16'hFEC3;    16'd12275: out <= 16'h040F;
    16'd12276: out <= 16'h01C6;    16'd12277: out <= 16'h02BA;    16'd12278: out <= 16'hFFC1;    16'd12279: out <= 16'hFA49;
    16'd12280: out <= 16'hFF26;    16'd12281: out <= 16'hFC15;    16'd12282: out <= 16'h0842;    16'd12283: out <= 16'hFFDC;
    16'd12284: out <= 16'hFF9E;    16'd12285: out <= 16'h01BE;    16'd12286: out <= 16'hF978;    16'd12287: out <= 16'h0443;
    16'd12288: out <= 16'hFE56;    16'd12289: out <= 16'h0115;    16'd12290: out <= 16'h08FF;    16'd12291: out <= 16'h02A5;
    16'd12292: out <= 16'h00E3;    16'd12293: out <= 16'hFAC7;    16'd12294: out <= 16'hFC38;    16'd12295: out <= 16'h021C;
    16'd12296: out <= 16'hFE62;    16'd12297: out <= 16'h0235;    16'd12298: out <= 16'hF856;    16'd12299: out <= 16'hFF41;
    16'd12300: out <= 16'hFD53;    16'd12301: out <= 16'hFE7D;    16'd12302: out <= 16'h0348;    16'd12303: out <= 16'hFD19;
    16'd12304: out <= 16'hFD1F;    16'd12305: out <= 16'h019E;    16'd12306: out <= 16'h01D9;    16'd12307: out <= 16'h0187;
    16'd12308: out <= 16'h0048;    16'd12309: out <= 16'hFF46;    16'd12310: out <= 16'h0157;    16'd12311: out <= 16'hFF5D;
    16'd12312: out <= 16'hF9E1;    16'd12313: out <= 16'h0295;    16'd12314: out <= 16'h03E0;    16'd12315: out <= 16'hFC9F;
    16'd12316: out <= 16'h00F6;    16'd12317: out <= 16'h086C;    16'd12318: out <= 16'h01A1;    16'd12319: out <= 16'h024D;
    16'd12320: out <= 16'hFDB1;    16'd12321: out <= 16'hFDC0;    16'd12322: out <= 16'h038F;    16'd12323: out <= 16'h0349;
    16'd12324: out <= 16'h02D5;    16'd12325: out <= 16'h0024;    16'd12326: out <= 16'h023B;    16'd12327: out <= 16'h074D;
    16'd12328: out <= 16'h025B;    16'd12329: out <= 16'h0471;    16'd12330: out <= 16'h06A1;    16'd12331: out <= 16'h0325;
    16'd12332: out <= 16'h062B;    16'd12333: out <= 16'h0503;    16'd12334: out <= 16'h00CB;    16'd12335: out <= 16'h01ED;
    16'd12336: out <= 16'h02B5;    16'd12337: out <= 16'h006D;    16'd12338: out <= 16'h02E7;    16'd12339: out <= 16'h00EA;
    16'd12340: out <= 16'h0516;    16'd12341: out <= 16'h06CB;    16'd12342: out <= 16'h04FE;    16'd12343: out <= 16'h03D5;
    16'd12344: out <= 16'h049B;    16'd12345: out <= 16'h065E;    16'd12346: out <= 16'h023E;    16'd12347: out <= 16'h07BC;
    16'd12348: out <= 16'hFFDC;    16'd12349: out <= 16'h0470;    16'd12350: out <= 16'h046C;    16'd12351: out <= 16'h05C3;
    16'd12352: out <= 16'h03FB;    16'd12353: out <= 16'h0534;    16'd12354: out <= 16'h064D;    16'd12355: out <= 16'h070C;
    16'd12356: out <= 16'h0069;    16'd12357: out <= 16'h027A;    16'd12358: out <= 16'h024A;    16'd12359: out <= 16'h0B08;
    16'd12360: out <= 16'h0152;    16'd12361: out <= 16'h03B7;    16'd12362: out <= 16'h00A5;    16'd12363: out <= 16'h0199;
    16'd12364: out <= 16'h04BC;    16'd12365: out <= 16'h00CC;    16'd12366: out <= 16'hFEF4;    16'd12367: out <= 16'h021F;
    16'd12368: out <= 16'h01A5;    16'd12369: out <= 16'h0B17;    16'd12370: out <= 16'h048B;    16'd12371: out <= 16'h02E3;
    16'd12372: out <= 16'h0921;    16'd12373: out <= 16'hFF93;    16'd12374: out <= 16'h06FF;    16'd12375: out <= 16'h037B;
    16'd12376: out <= 16'h00E4;    16'd12377: out <= 16'h0C09;    16'd12378: out <= 16'h01D0;    16'd12379: out <= 16'h02EA;
    16'd12380: out <= 16'hFF32;    16'd12381: out <= 16'h0ABF;    16'd12382: out <= 16'h07C5;    16'd12383: out <= 16'h0617;
    16'd12384: out <= 16'h06A5;    16'd12385: out <= 16'h0321;    16'd12386: out <= 16'h017D;    16'd12387: out <= 16'hFDDC;
    16'd12388: out <= 16'hFE3E;    16'd12389: out <= 16'hFF1D;    16'd12390: out <= 16'hFFCF;    16'd12391: out <= 16'h0457;
    16'd12392: out <= 16'h021B;    16'd12393: out <= 16'h098A;    16'd12394: out <= 16'hFB82;    16'd12395: out <= 16'hFF2D;
    16'd12396: out <= 16'hFBEF;    16'd12397: out <= 16'h05B2;    16'd12398: out <= 16'hF98B;    16'd12399: out <= 16'h0158;
    16'd12400: out <= 16'h03FA;    16'd12401: out <= 16'h0605;    16'd12402: out <= 16'h040A;    16'd12403: out <= 16'hFD91;
    16'd12404: out <= 16'h0500;    16'd12405: out <= 16'h06F0;    16'd12406: out <= 16'h0010;    16'd12407: out <= 16'h0364;
    16'd12408: out <= 16'h03BA;    16'd12409: out <= 16'h0477;    16'd12410: out <= 16'h002B;    16'd12411: out <= 16'hFF69;
    16'd12412: out <= 16'h0548;    16'd12413: out <= 16'h02FE;    16'd12414: out <= 16'h098B;    16'd12415: out <= 16'h0DA2;
    16'd12416: out <= 16'h059B;    16'd12417: out <= 16'h0607;    16'd12418: out <= 16'h026D;    16'd12419: out <= 16'h0273;
    16'd12420: out <= 16'h0A59;    16'd12421: out <= 16'hFCE3;    16'd12422: out <= 16'hFFDF;    16'd12423: out <= 16'h0A33;
    16'd12424: out <= 16'h0155;    16'd12425: out <= 16'h041D;    16'd12426: out <= 16'h0910;    16'd12427: out <= 16'h023E;
    16'd12428: out <= 16'h0699;    16'd12429: out <= 16'h0376;    16'd12430: out <= 16'h016A;    16'd12431: out <= 16'hFE75;
    16'd12432: out <= 16'h03BA;    16'd12433: out <= 16'h06F9;    16'd12434: out <= 16'h07C7;    16'd12435: out <= 16'h05EF;
    16'd12436: out <= 16'hFF05;    16'd12437: out <= 16'h04C8;    16'd12438: out <= 16'h00E6;    16'd12439: out <= 16'h00C8;
    16'd12440: out <= 16'hFE04;    16'd12441: out <= 16'h07EB;    16'd12442: out <= 16'h0000;    16'd12443: out <= 16'hFEA0;
    16'd12444: out <= 16'h0425;    16'd12445: out <= 16'h00DC;    16'd12446: out <= 16'h06E6;    16'd12447: out <= 16'hFE29;
    16'd12448: out <= 16'h0278;    16'd12449: out <= 16'hFE7C;    16'd12450: out <= 16'h0049;    16'd12451: out <= 16'h01D3;
    16'd12452: out <= 16'h05D9;    16'd12453: out <= 16'h0151;    16'd12454: out <= 16'h0578;    16'd12455: out <= 16'h08D5;
    16'd12456: out <= 16'h03F2;    16'd12457: out <= 16'h0411;    16'd12458: out <= 16'h020F;    16'd12459: out <= 16'h099E;
    16'd12460: out <= 16'h02D0;    16'd12461: out <= 16'h067F;    16'd12462: out <= 16'h0263;    16'd12463: out <= 16'h07FF;
    16'd12464: out <= 16'h0351;    16'd12465: out <= 16'h02B9;    16'd12466: out <= 16'h01D4;    16'd12467: out <= 16'h0551;
    16'd12468: out <= 16'h0251;    16'd12469: out <= 16'h0A65;    16'd12470: out <= 16'h03DF;    16'd12471: out <= 16'h07C1;
    16'd12472: out <= 16'h04E8;    16'd12473: out <= 16'hFF50;    16'd12474: out <= 16'h01C8;    16'd12475: out <= 16'h09D4;
    16'd12476: out <= 16'h05C5;    16'd12477: out <= 16'hFF3B;    16'd12478: out <= 16'h09FD;    16'd12479: out <= 16'h050E;
    16'd12480: out <= 16'h01D1;    16'd12481: out <= 16'h03C9;    16'd12482: out <= 16'h0897;    16'd12483: out <= 16'hFF16;
    16'd12484: out <= 16'h0930;    16'd12485: out <= 16'h03B9;    16'd12486: out <= 16'h070B;    16'd12487: out <= 16'h0995;
    16'd12488: out <= 16'h06E2;    16'd12489: out <= 16'h06CD;    16'd12490: out <= 16'h0C04;    16'd12491: out <= 16'h0894;
    16'd12492: out <= 16'h0461;    16'd12493: out <= 16'h079B;    16'd12494: out <= 16'h03AE;    16'd12495: out <= 16'h07CD;
    16'd12496: out <= 16'h01C3;    16'd12497: out <= 16'h0607;    16'd12498: out <= 16'hFD01;    16'd12499: out <= 16'h0AD3;
    16'd12500: out <= 16'h02F6;    16'd12501: out <= 16'h021D;    16'd12502: out <= 16'h0439;    16'd12503: out <= 16'h050B;
    16'd12504: out <= 16'h01DB;    16'd12505: out <= 16'hFCED;    16'd12506: out <= 16'hF85B;    16'd12507: out <= 16'h01E8;
    16'd12508: out <= 16'hFCF9;    16'd12509: out <= 16'hFF57;    16'd12510: out <= 16'h028A;    16'd12511: out <= 16'h02D6;
    16'd12512: out <= 16'h01E1;    16'd12513: out <= 16'h005F;    16'd12514: out <= 16'h093F;    16'd12515: out <= 16'hFC09;
    16'd12516: out <= 16'h0521;    16'd12517: out <= 16'hF997;    16'd12518: out <= 16'hF7E5;    16'd12519: out <= 16'hFB46;
    16'd12520: out <= 16'h0735;    16'd12521: out <= 16'hFE05;    16'd12522: out <= 16'hF9D0;    16'd12523: out <= 16'h0116;
    16'd12524: out <= 16'h01ED;    16'd12525: out <= 16'hFCCC;    16'd12526: out <= 16'hFCD2;    16'd12527: out <= 16'hFF6A;
    16'd12528: out <= 16'h023D;    16'd12529: out <= 16'hFE81;    16'd12530: out <= 16'hF8CE;    16'd12531: out <= 16'h00A8;
    16'd12532: out <= 16'h0017;    16'd12533: out <= 16'h0386;    16'd12534: out <= 16'h0D55;    16'd12535: out <= 16'hFA69;
    16'd12536: out <= 16'h053C;    16'd12537: out <= 16'h059C;    16'd12538: out <= 16'h0AA3;    16'd12539: out <= 16'hFEDE;
    16'd12540: out <= 16'h0112;    16'd12541: out <= 16'h0141;    16'd12542: out <= 16'h0128;    16'd12543: out <= 16'h0426;
    16'd12544: out <= 16'hFBD7;    16'd12545: out <= 16'hFD88;    16'd12546: out <= 16'h040F;    16'd12547: out <= 16'h0397;
    16'd12548: out <= 16'h0342;    16'd12549: out <= 16'hFC32;    16'd12550: out <= 16'h0075;    16'd12551: out <= 16'hFBF3;
    16'd12552: out <= 16'h01E7;    16'd12553: out <= 16'h037C;    16'd12554: out <= 16'hFE17;    16'd12555: out <= 16'h045B;
    16'd12556: out <= 16'h023E;    16'd12557: out <= 16'hFCB1;    16'd12558: out <= 16'hFF65;    16'd12559: out <= 16'h00C0;
    16'd12560: out <= 16'hFEC2;    16'd12561: out <= 16'h067E;    16'd12562: out <= 16'h0111;    16'd12563: out <= 16'h009F;
    16'd12564: out <= 16'hFCF3;    16'd12565: out <= 16'h079E;    16'd12566: out <= 16'h054B;    16'd12567: out <= 16'h00BB;
    16'd12568: out <= 16'hFC9F;    16'd12569: out <= 16'hFFB2;    16'd12570: out <= 16'h02E1;    16'd12571: out <= 16'h05E1;
    16'd12572: out <= 16'hFD4C;    16'd12573: out <= 16'h02F1;    16'd12574: out <= 16'h0328;    16'd12575: out <= 16'hFDFF;
    16'd12576: out <= 16'h01A9;    16'd12577: out <= 16'hFE9D;    16'd12578: out <= 16'h0254;    16'd12579: out <= 16'h05EA;
    16'd12580: out <= 16'hFD3F;    16'd12581: out <= 16'h044E;    16'd12582: out <= 16'h0509;    16'd12583: out <= 16'h011E;
    16'd12584: out <= 16'h044B;    16'd12585: out <= 16'hFE96;    16'd12586: out <= 16'h089E;    16'd12587: out <= 16'h0CB3;
    16'd12588: out <= 16'h04CB;    16'd12589: out <= 16'h0BF0;    16'd12590: out <= 16'hFD07;    16'd12591: out <= 16'h06C1;
    16'd12592: out <= 16'h01FE;    16'd12593: out <= 16'h082F;    16'd12594: out <= 16'h0808;    16'd12595: out <= 16'hFD2E;
    16'd12596: out <= 16'h063D;    16'd12597: out <= 16'h0070;    16'd12598: out <= 16'h0382;    16'd12599: out <= 16'h0532;
    16'd12600: out <= 16'h0266;    16'd12601: out <= 16'h0209;    16'd12602: out <= 16'h07B2;    16'd12603: out <= 16'h034A;
    16'd12604: out <= 16'h01AE;    16'd12605: out <= 16'h0446;    16'd12606: out <= 16'h0721;    16'd12607: out <= 16'h0276;
    16'd12608: out <= 16'h038F;    16'd12609: out <= 16'h021C;    16'd12610: out <= 16'h0365;    16'd12611: out <= 16'h03ED;
    16'd12612: out <= 16'hF9E1;    16'd12613: out <= 16'h02DC;    16'd12614: out <= 16'h01F4;    16'd12615: out <= 16'h08A7;
    16'd12616: out <= 16'h012F;    16'd12617: out <= 16'hFEF8;    16'd12618: out <= 16'h01C4;    16'd12619: out <= 16'h059D;
    16'd12620: out <= 16'h0806;    16'd12621: out <= 16'h027F;    16'd12622: out <= 16'hFDC0;    16'd12623: out <= 16'h0066;
    16'd12624: out <= 16'h02E3;    16'd12625: out <= 16'hFFE1;    16'd12626: out <= 16'h0301;    16'd12627: out <= 16'h0D8A;
    16'd12628: out <= 16'h0474;    16'd12629: out <= 16'h0C20;    16'd12630: out <= 16'hFE63;    16'd12631: out <= 16'hFB1F;
    16'd12632: out <= 16'h035D;    16'd12633: out <= 16'h0109;    16'd12634: out <= 16'h0694;    16'd12635: out <= 16'h02AA;
    16'd12636: out <= 16'hFF7D;    16'd12637: out <= 16'hFD3C;    16'd12638: out <= 16'h04F7;    16'd12639: out <= 16'hFFA4;
    16'd12640: out <= 16'h08B5;    16'd12641: out <= 16'hFDF4;    16'd12642: out <= 16'hFD31;    16'd12643: out <= 16'hFF7F;
    16'd12644: out <= 16'hFE2C;    16'd12645: out <= 16'h0691;    16'd12646: out <= 16'h0571;    16'd12647: out <= 16'hFFCD;
    16'd12648: out <= 16'h00BC;    16'd12649: out <= 16'h051F;    16'd12650: out <= 16'hFE93;    16'd12651: out <= 16'hFFED;
    16'd12652: out <= 16'h0411;    16'd12653: out <= 16'h0011;    16'd12654: out <= 16'h04B8;    16'd12655: out <= 16'h0464;
    16'd12656: out <= 16'h043D;    16'd12657: out <= 16'h0177;    16'd12658: out <= 16'h02D8;    16'd12659: out <= 16'h026C;
    16'd12660: out <= 16'h04D9;    16'd12661: out <= 16'h05EA;    16'd12662: out <= 16'h0837;    16'd12663: out <= 16'hFF1A;
    16'd12664: out <= 16'h0893;    16'd12665: out <= 16'h084E;    16'd12666: out <= 16'h0302;    16'd12667: out <= 16'h08E5;
    16'd12668: out <= 16'hFEEA;    16'd12669: out <= 16'h07DA;    16'd12670: out <= 16'h0529;    16'd12671: out <= 16'h096F;
    16'd12672: out <= 16'h0293;    16'd12673: out <= 16'h00E6;    16'd12674: out <= 16'hFF4E;    16'd12675: out <= 16'hFF69;
    16'd12676: out <= 16'h09FA;    16'd12677: out <= 16'h03C5;    16'd12678: out <= 16'h029B;    16'd12679: out <= 16'h0441;
    16'd12680: out <= 16'h0C11;    16'd12681: out <= 16'hFFF7;    16'd12682: out <= 16'hFC48;    16'd12683: out <= 16'h016B;
    16'd12684: out <= 16'h09EC;    16'd12685: out <= 16'hFDA6;    16'd12686: out <= 16'h0563;    16'd12687: out <= 16'hFDD3;
    16'd12688: out <= 16'h0594;    16'd12689: out <= 16'h072F;    16'd12690: out <= 16'h0C56;    16'd12691: out <= 16'h0667;
    16'd12692: out <= 16'h029E;    16'd12693: out <= 16'h045B;    16'd12694: out <= 16'h023D;    16'd12695: out <= 16'h03EB;
    16'd12696: out <= 16'h02E6;    16'd12697: out <= 16'h067D;    16'd12698: out <= 16'h02F5;    16'd12699: out <= 16'h023F;
    16'd12700: out <= 16'hFFDD;    16'd12701: out <= 16'h0675;    16'd12702: out <= 16'h0709;    16'd12703: out <= 16'h0117;
    16'd12704: out <= 16'h0670;    16'd12705: out <= 16'h06FD;    16'd12706: out <= 16'h02B8;    16'd12707: out <= 16'h0185;
    16'd12708: out <= 16'hFF72;    16'd12709: out <= 16'h068B;    16'd12710: out <= 16'hFD7F;    16'd12711: out <= 16'h08BF;
    16'd12712: out <= 16'h079A;    16'd12713: out <= 16'h065F;    16'd12714: out <= 16'h03A8;    16'd12715: out <= 16'h0258;
    16'd12716: out <= 16'h0394;    16'd12717: out <= 16'hFDB2;    16'd12718: out <= 16'h02CB;    16'd12719: out <= 16'h08D1;
    16'd12720: out <= 16'h063A;    16'd12721: out <= 16'h08A8;    16'd12722: out <= 16'hFF5A;    16'd12723: out <= 16'h0325;
    16'd12724: out <= 16'h069A;    16'd12725: out <= 16'h0454;    16'd12726: out <= 16'hFF94;    16'd12727: out <= 16'hFDEC;
    16'd12728: out <= 16'hFE0D;    16'd12729: out <= 16'hFF96;    16'd12730: out <= 16'h04FF;    16'd12731: out <= 16'h03FB;
    16'd12732: out <= 16'h0607;    16'd12733: out <= 16'h084F;    16'd12734: out <= 16'h0216;    16'd12735: out <= 16'h020A;
    16'd12736: out <= 16'h0832;    16'd12737: out <= 16'h02E9;    16'd12738: out <= 16'h01FE;    16'd12739: out <= 16'h0072;
    16'd12740: out <= 16'h02F6;    16'd12741: out <= 16'h048B;    16'd12742: out <= 16'hFB78;    16'd12743: out <= 16'h0308;
    16'd12744: out <= 16'h0433;    16'd12745: out <= 16'h07BB;    16'd12746: out <= 16'h0083;    16'd12747: out <= 16'h04FA;
    16'd12748: out <= 16'h0471;    16'd12749: out <= 16'h01D7;    16'd12750: out <= 16'h02D8;    16'd12751: out <= 16'h050E;
    16'd12752: out <= 16'h0135;    16'd12753: out <= 16'hFBBA;    16'd12754: out <= 16'h0C1A;    16'd12755: out <= 16'h0312;
    16'd12756: out <= 16'hFEE2;    16'd12757: out <= 16'h0602;    16'd12758: out <= 16'h0441;    16'd12759: out <= 16'h04B6;
    16'd12760: out <= 16'h079A;    16'd12761: out <= 16'h0095;    16'd12762: out <= 16'hFD04;    16'd12763: out <= 16'h01F1;
    16'd12764: out <= 16'hFFA3;    16'd12765: out <= 16'h00AB;    16'd12766: out <= 16'hFF45;    16'd12767: out <= 16'hFF44;
    16'd12768: out <= 16'hFDAE;    16'd12769: out <= 16'hFAE4;    16'd12770: out <= 16'hF925;    16'd12771: out <= 16'h0615;
    16'd12772: out <= 16'h031B;    16'd12773: out <= 16'hFBE6;    16'd12774: out <= 16'hFCE1;    16'd12775: out <= 16'hFC98;
    16'd12776: out <= 16'hFE48;    16'd12777: out <= 16'h02AA;    16'd12778: out <= 16'hFCE9;    16'd12779: out <= 16'h03C0;
    16'd12780: out <= 16'hFF5C;    16'd12781: out <= 16'h013E;    16'd12782: out <= 16'h0796;    16'd12783: out <= 16'hFEB0;
    16'd12784: out <= 16'hFEC7;    16'd12785: out <= 16'hFB58;    16'd12786: out <= 16'hFBD6;    16'd12787: out <= 16'hFA01;
    16'd12788: out <= 16'hFB28;    16'd12789: out <= 16'h027A;    16'd12790: out <= 16'hFEF3;    16'd12791: out <= 16'h07A9;
    16'd12792: out <= 16'h0198;    16'd12793: out <= 16'hF83D;    16'd12794: out <= 16'h02A9;    16'd12795: out <= 16'hFFFD;
    16'd12796: out <= 16'h03BB;    16'd12797: out <= 16'hFF95;    16'd12798: out <= 16'h0667;    16'd12799: out <= 16'hFDAC;
    16'd12800: out <= 16'hFABF;    16'd12801: out <= 16'h04F8;    16'd12802: out <= 16'h010A;    16'd12803: out <= 16'h07E7;
    16'd12804: out <= 16'hFB23;    16'd12805: out <= 16'h058E;    16'd12806: out <= 16'h0445;    16'd12807: out <= 16'h02FE;
    16'd12808: out <= 16'h01E1;    16'd12809: out <= 16'hFFC9;    16'd12810: out <= 16'h002B;    16'd12811: out <= 16'hFC1D;
    16'd12812: out <= 16'h06BA;    16'd12813: out <= 16'h061E;    16'd12814: out <= 16'h0433;    16'd12815: out <= 16'hFFA9;
    16'd12816: out <= 16'hFDF4;    16'd12817: out <= 16'hFE6A;    16'd12818: out <= 16'h0242;    16'd12819: out <= 16'h04E5;
    16'd12820: out <= 16'hFDCF;    16'd12821: out <= 16'hFF9C;    16'd12822: out <= 16'h0706;    16'd12823: out <= 16'hFB9A;
    16'd12824: out <= 16'h009E;    16'd12825: out <= 16'hFD24;    16'd12826: out <= 16'h0280;    16'd12827: out <= 16'hFEFB;
    16'd12828: out <= 16'h03EF;    16'd12829: out <= 16'hFF59;    16'd12830: out <= 16'h001F;    16'd12831: out <= 16'h04E7;
    16'd12832: out <= 16'hFF4B;    16'd12833: out <= 16'h0208;    16'd12834: out <= 16'hFCC9;    16'd12835: out <= 16'hFA71;
    16'd12836: out <= 16'hF821;    16'd12837: out <= 16'h0197;    16'd12838: out <= 16'hFC96;    16'd12839: out <= 16'h0627;
    16'd12840: out <= 16'h053B;    16'd12841: out <= 16'h0104;    16'd12842: out <= 16'hFC39;    16'd12843: out <= 16'h033B;
    16'd12844: out <= 16'h05BD;    16'd12845: out <= 16'h04C1;    16'd12846: out <= 16'h01FF;    16'd12847: out <= 16'h07DC;
    16'd12848: out <= 16'h0343;    16'd12849: out <= 16'h0943;    16'd12850: out <= 16'h04F8;    16'd12851: out <= 16'h07BE;
    16'd12852: out <= 16'h0341;    16'd12853: out <= 16'h0B3B;    16'd12854: out <= 16'h0306;    16'd12855: out <= 16'h0566;
    16'd12856: out <= 16'hFEF9;    16'd12857: out <= 16'h0310;    16'd12858: out <= 16'h0724;    16'd12859: out <= 16'h07CD;
    16'd12860: out <= 16'h078D;    16'd12861: out <= 16'h06D5;    16'd12862: out <= 16'hFF55;    16'd12863: out <= 16'h0A8F;
    16'd12864: out <= 16'h0C33;    16'd12865: out <= 16'hFFA3;    16'd12866: out <= 16'h0739;    16'd12867: out <= 16'h07FF;
    16'd12868: out <= 16'h00AD;    16'd12869: out <= 16'hFE1A;    16'd12870: out <= 16'h0B7A;    16'd12871: out <= 16'h02C6;
    16'd12872: out <= 16'h0C11;    16'd12873: out <= 16'h0766;    16'd12874: out <= 16'h02C5;    16'd12875: out <= 16'h08A6;
    16'd12876: out <= 16'h0630;    16'd12877: out <= 16'h0776;    16'd12878: out <= 16'h016B;    16'd12879: out <= 16'h0C21;
    16'd12880: out <= 16'hFF4E;    16'd12881: out <= 16'h07F4;    16'd12882: out <= 16'h0798;    16'd12883: out <= 16'hFD7E;
    16'd12884: out <= 16'hFD75;    16'd12885: out <= 16'h048F;    16'd12886: out <= 16'h08E7;    16'd12887: out <= 16'hFE91;
    16'd12888: out <= 16'h0B43;    16'd12889: out <= 16'h0509;    16'd12890: out <= 16'h0507;    16'd12891: out <= 16'h0888;
    16'd12892: out <= 16'h0272;    16'd12893: out <= 16'h04AA;    16'd12894: out <= 16'hFE9D;    16'd12895: out <= 16'h0022;
    16'd12896: out <= 16'h0050;    16'd12897: out <= 16'h0571;    16'd12898: out <= 16'h031D;    16'd12899: out <= 16'hF903;
    16'd12900: out <= 16'h02CF;    16'd12901: out <= 16'h03E4;    16'd12902: out <= 16'h0AEF;    16'd12903: out <= 16'hFDB0;
    16'd12904: out <= 16'h02AD;    16'd12905: out <= 16'h0796;    16'd12906: out <= 16'h049A;    16'd12907: out <= 16'h0195;
    16'd12908: out <= 16'hFD04;    16'd12909: out <= 16'h071F;    16'd12910: out <= 16'h053F;    16'd12911: out <= 16'h05A1;
    16'd12912: out <= 16'h00B3;    16'd12913: out <= 16'hFFED;    16'd12914: out <= 16'h0493;    16'd12915: out <= 16'h02AE;
    16'd12916: out <= 16'h00FB;    16'd12917: out <= 16'h0769;    16'd12918: out <= 16'h0273;    16'd12919: out <= 16'h0365;
    16'd12920: out <= 16'h024E;    16'd12921: out <= 16'h0423;    16'd12922: out <= 16'h03A9;    16'd12923: out <= 16'h0491;
    16'd12924: out <= 16'h0D98;    16'd12925: out <= 16'h0440;    16'd12926: out <= 16'h0501;    16'd12927: out <= 16'h0AF4;
    16'd12928: out <= 16'h0A49;    16'd12929: out <= 16'h04B4;    16'd12930: out <= 16'h0259;    16'd12931: out <= 16'h02E6;
    16'd12932: out <= 16'h02E3;    16'd12933: out <= 16'h06EA;    16'd12934: out <= 16'h0515;    16'd12935: out <= 16'hFFD8;
    16'd12936: out <= 16'h05D9;    16'd12937: out <= 16'h0425;    16'd12938: out <= 16'h04FD;    16'd12939: out <= 16'h02DF;
    16'd12940: out <= 16'h027E;    16'd12941: out <= 16'h00FF;    16'd12942: out <= 16'h0102;    16'd12943: out <= 16'h0B8C;
    16'd12944: out <= 16'h00AC;    16'd12945: out <= 16'h0230;    16'd12946: out <= 16'h051D;    16'd12947: out <= 16'h026A;
    16'd12948: out <= 16'h0290;    16'd12949: out <= 16'h01C5;    16'd12950: out <= 16'h054D;    16'd12951: out <= 16'h05DB;
    16'd12952: out <= 16'h07A7;    16'd12953: out <= 16'hFF77;    16'd12954: out <= 16'hFECB;    16'd12955: out <= 16'h00DA;
    16'd12956: out <= 16'h08E1;    16'd12957: out <= 16'h0991;    16'd12958: out <= 16'h0300;    16'd12959: out <= 16'hFF87;
    16'd12960: out <= 16'hFF78;    16'd12961: out <= 16'hFCBA;    16'd12962: out <= 16'h0616;    16'd12963: out <= 16'h067F;
    16'd12964: out <= 16'h05FE;    16'd12965: out <= 16'h0911;    16'd12966: out <= 16'h03B9;    16'd12967: out <= 16'h04F8;
    16'd12968: out <= 16'hFBDC;    16'd12969: out <= 16'hFE4E;    16'd12970: out <= 16'hFDB6;    16'd12971: out <= 16'hFD5E;
    16'd12972: out <= 16'h0311;    16'd12973: out <= 16'h055E;    16'd12974: out <= 16'h0351;    16'd12975: out <= 16'h0702;
    16'd12976: out <= 16'h040B;    16'd12977: out <= 16'h0636;    16'd12978: out <= 16'hF47D;    16'd12979: out <= 16'h071A;
    16'd12980: out <= 16'h07A6;    16'd12981: out <= 16'h0093;    16'd12982: out <= 16'h0562;    16'd12983: out <= 16'h0343;
    16'd12984: out <= 16'h0178;    16'd12985: out <= 16'h04D3;    16'd12986: out <= 16'h0343;    16'd12987: out <= 16'hFE93;
    16'd12988: out <= 16'h01A3;    16'd12989: out <= 16'h04C4;    16'd12990: out <= 16'h0238;    16'd12991: out <= 16'h074F;
    16'd12992: out <= 16'h0A66;    16'd12993: out <= 16'h01AA;    16'd12994: out <= 16'h0A67;    16'd12995: out <= 16'h0033;
    16'd12996: out <= 16'h026F;    16'd12997: out <= 16'hFD1C;    16'd12998: out <= 16'h00FB;    16'd12999: out <= 16'h0A2F;
    16'd13000: out <= 16'h0667;    16'd13001: out <= 16'h07F8;    16'd13002: out <= 16'h0632;    16'd13003: out <= 16'h083A;
    16'd13004: out <= 16'h061A;    16'd13005: out <= 16'h0196;    16'd13006: out <= 16'hFF56;    16'd13007: out <= 16'h03DA;
    16'd13008: out <= 16'h03CF;    16'd13009: out <= 16'h02F4;    16'd13010: out <= 16'h030E;    16'd13011: out <= 16'h05F8;
    16'd13012: out <= 16'h023B;    16'd13013: out <= 16'hFD74;    16'd13014: out <= 16'h05D0;    16'd13015: out <= 16'hFFC4;
    16'd13016: out <= 16'hFCAC;    16'd13017: out <= 16'hFFD1;    16'd13018: out <= 16'h0729;    16'd13019: out <= 16'h08D0;
    16'd13020: out <= 16'hFBD5;    16'd13021: out <= 16'h079F;    16'd13022: out <= 16'hFF76;    16'd13023: out <= 16'h0404;
    16'd13024: out <= 16'hFF4A;    16'd13025: out <= 16'hFC0E;    16'd13026: out <= 16'h007A;    16'd13027: out <= 16'hFF81;
    16'd13028: out <= 16'hFE2E;    16'd13029: out <= 16'h001E;    16'd13030: out <= 16'h004E;    16'd13031: out <= 16'h0119;
    16'd13032: out <= 16'h001E;    16'd13033: out <= 16'hFBE6;    16'd13034: out <= 16'h01A7;    16'd13035: out <= 16'hFF1C;
    16'd13036: out <= 16'hFE70;    16'd13037: out <= 16'hFF12;    16'd13038: out <= 16'hFBE3;    16'd13039: out <= 16'hFE77;
    16'd13040: out <= 16'hF753;    16'd13041: out <= 16'h0456;    16'd13042: out <= 16'hFD0D;    16'd13043: out <= 16'hFEE0;
    16'd13044: out <= 16'h00C9;    16'd13045: out <= 16'h078E;    16'd13046: out <= 16'h0A7E;    16'd13047: out <= 16'hFA55;
    16'd13048: out <= 16'hFD55;    16'd13049: out <= 16'hFC0B;    16'd13050: out <= 16'h051C;    16'd13051: out <= 16'hFCFF;
    16'd13052: out <= 16'hFCBF;    16'd13053: out <= 16'h05FE;    16'd13054: out <= 16'h0067;    16'd13055: out <= 16'hF7A8;
    16'd13056: out <= 16'h00CD;    16'd13057: out <= 16'hFF93;    16'd13058: out <= 16'h03D6;    16'd13059: out <= 16'hFA09;
    16'd13060: out <= 16'h04B7;    16'd13061: out <= 16'h0174;    16'd13062: out <= 16'hFFED;    16'd13063: out <= 16'h030E;
    16'd13064: out <= 16'hFEAA;    16'd13065: out <= 16'h01F4;    16'd13066: out <= 16'hFB1C;    16'd13067: out <= 16'h019F;
    16'd13068: out <= 16'h04DD;    16'd13069: out <= 16'h0516;    16'd13070: out <= 16'h0284;    16'd13071: out <= 16'h0380;
    16'd13072: out <= 16'hFF1C;    16'd13073: out <= 16'h0424;    16'd13074: out <= 16'h04C3;    16'd13075: out <= 16'h04B2;
    16'd13076: out <= 16'h01FD;    16'd13077: out <= 16'h0751;    16'd13078: out <= 16'hF7D0;    16'd13079: out <= 16'hFBC4;
    16'd13080: out <= 16'h0125;    16'd13081: out <= 16'h0223;    16'd13082: out <= 16'hFC9B;    16'd13083: out <= 16'hFFAE;
    16'd13084: out <= 16'hFD8D;    16'd13085: out <= 16'hFD4D;    16'd13086: out <= 16'hFF64;    16'd13087: out <= 16'h01E1;
    16'd13088: out <= 16'h027B;    16'd13089: out <= 16'hFED3;    16'd13090: out <= 16'h0076;    16'd13091: out <= 16'h0331;
    16'd13092: out <= 16'hF6AD;    16'd13093: out <= 16'hFE34;    16'd13094: out <= 16'h02B5;    16'd13095: out <= 16'h0A24;
    16'd13096: out <= 16'h08A9;    16'd13097: out <= 16'h026B;    16'd13098: out <= 16'h02BD;    16'd13099: out <= 16'h010E;
    16'd13100: out <= 16'h01A6;    16'd13101: out <= 16'h007D;    16'd13102: out <= 16'h04FA;    16'd13103: out <= 16'h0070;
    16'd13104: out <= 16'hFEB9;    16'd13105: out <= 16'h0A92;    16'd13106: out <= 16'h0439;    16'd13107: out <= 16'hF9BD;
    16'd13108: out <= 16'hF9B8;    16'd13109: out <= 16'h05BF;    16'd13110: out <= 16'h026F;    16'd13111: out <= 16'h0667;
    16'd13112: out <= 16'h03BA;    16'd13113: out <= 16'h07DF;    16'd13114: out <= 16'hFFBC;    16'd13115: out <= 16'h002F;
    16'd13116: out <= 16'h0288;    16'd13117: out <= 16'hF7F0;    16'd13118: out <= 16'h03EC;    16'd13119: out <= 16'h01CC;
    16'd13120: out <= 16'h0117;    16'd13121: out <= 16'h0202;    16'd13122: out <= 16'h071E;    16'd13123: out <= 16'h0672;
    16'd13124: out <= 16'h03FD;    16'd13125: out <= 16'h059B;    16'd13126: out <= 16'h0273;    16'd13127: out <= 16'h01D1;
    16'd13128: out <= 16'h0095;    16'd13129: out <= 16'h0759;    16'd13130: out <= 16'hFEAD;    16'd13131: out <= 16'hFF8F;
    16'd13132: out <= 16'h06AA;    16'd13133: out <= 16'h0141;    16'd13134: out <= 16'h07C0;    16'd13135: out <= 16'h02DB;
    16'd13136: out <= 16'h098A;    16'd13137: out <= 16'h0448;    16'd13138: out <= 16'h0658;    16'd13139: out <= 16'h0C4D;
    16'd13140: out <= 16'h0A30;    16'd13141: out <= 16'h027D;    16'd13142: out <= 16'h0007;    16'd13143: out <= 16'h07C0;
    16'd13144: out <= 16'hFE46;    16'd13145: out <= 16'h10F5;    16'd13146: out <= 16'h0825;    16'd13147: out <= 16'h046D;
    16'd13148: out <= 16'hFF64;    16'd13149: out <= 16'hFD92;    16'd13150: out <= 16'h067D;    16'd13151: out <= 16'hFF2E;
    16'd13152: out <= 16'h0343;    16'd13153: out <= 16'h07ED;    16'd13154: out <= 16'h08EE;    16'd13155: out <= 16'h04AA;
    16'd13156: out <= 16'hFF2C;    16'd13157: out <= 16'h04E1;    16'd13158: out <= 16'h0255;    16'd13159: out <= 16'h08AC;
    16'd13160: out <= 16'h0249;    16'd13161: out <= 16'h064E;    16'd13162: out <= 16'h04BE;    16'd13163: out <= 16'h05B9;
    16'd13164: out <= 16'h0415;    16'd13165: out <= 16'h024D;    16'd13166: out <= 16'h0002;    16'd13167: out <= 16'h02A5;
    16'd13168: out <= 16'h056C;    16'd13169: out <= 16'h0853;    16'd13170: out <= 16'h02BD;    16'd13171: out <= 16'h09B1;
    16'd13172: out <= 16'hFFB0;    16'd13173: out <= 16'h0929;    16'd13174: out <= 16'h079C;    16'd13175: out <= 16'h09F3;
    16'd13176: out <= 16'h0387;    16'd13177: out <= 16'h0257;    16'd13178: out <= 16'h0387;    16'd13179: out <= 16'h016E;
    16'd13180: out <= 16'hFEF6;    16'd13181: out <= 16'h0302;    16'd13182: out <= 16'hFBC9;    16'd13183: out <= 16'h0712;
    16'd13184: out <= 16'h0562;    16'd13185: out <= 16'hFEF2;    16'd13186: out <= 16'h0412;    16'd13187: out <= 16'h00EE;
    16'd13188: out <= 16'h0270;    16'd13189: out <= 16'h0015;    16'd13190: out <= 16'h0807;    16'd13191: out <= 16'h05C6;
    16'd13192: out <= 16'h0421;    16'd13193: out <= 16'hFE8F;    16'd13194: out <= 16'h00A2;    16'd13195: out <= 16'h039D;
    16'd13196: out <= 16'h0477;    16'd13197: out <= 16'h0152;    16'd13198: out <= 16'h08D7;    16'd13199: out <= 16'h040F;
    16'd13200: out <= 16'h09CB;    16'd13201: out <= 16'h019F;    16'd13202: out <= 16'h0042;    16'd13203: out <= 16'hFE14;
    16'd13204: out <= 16'h0170;    16'd13205: out <= 16'h003B;    16'd13206: out <= 16'h0278;    16'd13207: out <= 16'hFE18;
    16'd13208: out <= 16'h0387;    16'd13209: out <= 16'h0877;    16'd13210: out <= 16'h0261;    16'd13211: out <= 16'h0664;
    16'd13212: out <= 16'h0BDA;    16'd13213: out <= 16'h0554;    16'd13214: out <= 16'h0A2C;    16'd13215: out <= 16'hFFBA;
    16'd13216: out <= 16'h04FB;    16'd13217: out <= 16'hFEF5;    16'd13218: out <= 16'h0242;    16'd13219: out <= 16'h080B;
    16'd13220: out <= 16'h07EB;    16'd13221: out <= 16'h00C3;    16'd13222: out <= 16'h0596;    16'd13223: out <= 16'h0769;
    16'd13224: out <= 16'h04B2;    16'd13225: out <= 16'h015A;    16'd13226: out <= 16'h09A5;    16'd13227: out <= 16'hFD5F;
    16'd13228: out <= 16'h052E;    16'd13229: out <= 16'h08E5;    16'd13230: out <= 16'h00A7;    16'd13231: out <= 16'h07DF;
    16'd13232: out <= 16'h095C;    16'd13233: out <= 16'h0308;    16'd13234: out <= 16'h02B2;    16'd13235: out <= 16'h0936;
    16'd13236: out <= 16'h018C;    16'd13237: out <= 16'hFE30;    16'd13238: out <= 16'h02D1;    16'd13239: out <= 16'h02F8;
    16'd13240: out <= 16'h01E2;    16'd13241: out <= 16'h0322;    16'd13242: out <= 16'h0276;    16'd13243: out <= 16'h078C;
    16'd13244: out <= 16'h03E2;    16'd13245: out <= 16'h036F;    16'd13246: out <= 16'hFB06;    16'd13247: out <= 16'h02F2;
    16'd13248: out <= 16'h05CE;    16'd13249: out <= 16'h04A1;    16'd13250: out <= 16'h0117;    16'd13251: out <= 16'h04D7;
    16'd13252: out <= 16'h06BA;    16'd13253: out <= 16'h0891;    16'd13254: out <= 16'hFF5D;    16'd13255: out <= 16'h0781;
    16'd13256: out <= 16'h0594;    16'd13257: out <= 16'h0260;    16'd13258: out <= 16'h005C;    16'd13259: out <= 16'h030D;
    16'd13260: out <= 16'h0099;    16'd13261: out <= 16'h04A1;    16'd13262: out <= 16'h0393;    16'd13263: out <= 16'h0654;
    16'd13264: out <= 16'hFDE4;    16'd13265: out <= 16'hFF5A;    16'd13266: out <= 16'h03E1;    16'd13267: out <= 16'hFFD9;
    16'd13268: out <= 16'h03BF;    16'd13269: out <= 16'hFF29;    16'd13270: out <= 16'h02DE;    16'd13271: out <= 16'h07A7;
    16'd13272: out <= 16'hFA50;    16'd13273: out <= 16'h0634;    16'd13274: out <= 16'h0165;    16'd13275: out <= 16'h052D;
    16'd13276: out <= 16'h0498;    16'd13277: out <= 16'hFE2E;    16'd13278: out <= 16'h0389;    16'd13279: out <= 16'h016B;
    16'd13280: out <= 16'hFD1C;    16'd13281: out <= 16'h0622;    16'd13282: out <= 16'h07A2;    16'd13283: out <= 16'hF3E2;
    16'd13284: out <= 16'hFF72;    16'd13285: out <= 16'h03B5;    16'd13286: out <= 16'hFEB0;    16'd13287: out <= 16'h03F7;
    16'd13288: out <= 16'hF5D6;    16'd13289: out <= 16'h0456;    16'd13290: out <= 16'hFE4B;    16'd13291: out <= 16'hFFFE;
    16'd13292: out <= 16'hF965;    16'd13293: out <= 16'hF8FB;    16'd13294: out <= 16'h0016;    16'd13295: out <= 16'h0205;
    16'd13296: out <= 16'h0437;    16'd13297: out <= 16'h04DA;    16'd13298: out <= 16'h0053;    16'd13299: out <= 16'h02C4;
    16'd13300: out <= 16'h06DE;    16'd13301: out <= 16'hFCDE;    16'd13302: out <= 16'hF9A8;    16'd13303: out <= 16'hFEC8;
    16'd13304: out <= 16'hFDDC;    16'd13305: out <= 16'hFF8B;    16'd13306: out <= 16'h02AE;    16'd13307: out <= 16'hFD69;
    16'd13308: out <= 16'h0718;    16'd13309: out <= 16'hFFBB;    16'd13310: out <= 16'hFFEE;    16'd13311: out <= 16'h033C;
    16'd13312: out <= 16'h039C;    16'd13313: out <= 16'hFD17;    16'd13314: out <= 16'hFFA0;    16'd13315: out <= 16'hFEA1;
    16'd13316: out <= 16'hFACF;    16'd13317: out <= 16'hFE57;    16'd13318: out <= 16'hFCEA;    16'd13319: out <= 16'hF8B3;
    16'd13320: out <= 16'h033C;    16'd13321: out <= 16'h0491;    16'd13322: out <= 16'hFF3E;    16'd13323: out <= 16'hFD35;
    16'd13324: out <= 16'h022B;    16'd13325: out <= 16'h00F7;    16'd13326: out <= 16'h0195;    16'd13327: out <= 16'h0787;
    16'd13328: out <= 16'h0252;    16'd13329: out <= 16'hFCBB;    16'd13330: out <= 16'hF9F0;    16'd13331: out <= 16'hFEA3;
    16'd13332: out <= 16'h02AC;    16'd13333: out <= 16'hFC98;    16'd13334: out <= 16'hFD6D;    16'd13335: out <= 16'hFA70;
    16'd13336: out <= 16'h0128;    16'd13337: out <= 16'h0177;    16'd13338: out <= 16'h0096;    16'd13339: out <= 16'hF9D1;
    16'd13340: out <= 16'hFB69;    16'd13341: out <= 16'hFB05;    16'd13342: out <= 16'h0397;    16'd13343: out <= 16'h010F;
    16'd13344: out <= 16'h05A3;    16'd13345: out <= 16'h06C9;    16'd13346: out <= 16'h0E09;    16'd13347: out <= 16'h0B56;
    16'd13348: out <= 16'hFC72;    16'd13349: out <= 16'hF9EF;    16'd13350: out <= 16'h049F;    16'd13351: out <= 16'h0575;
    16'd13352: out <= 16'h05D7;    16'd13353: out <= 16'h0688;    16'd13354: out <= 16'h055F;    16'd13355: out <= 16'h05A8;
    16'd13356: out <= 16'hFF63;    16'd13357: out <= 16'h0776;    16'd13358: out <= 16'h0420;    16'd13359: out <= 16'h041F;
    16'd13360: out <= 16'h069F;    16'd13361: out <= 16'h07A0;    16'd13362: out <= 16'h0642;    16'd13363: out <= 16'h0784;
    16'd13364: out <= 16'h00A2;    16'd13365: out <= 16'h0888;    16'd13366: out <= 16'h041D;    16'd13367: out <= 16'h0651;
    16'd13368: out <= 16'h0264;    16'd13369: out <= 16'h0292;    16'd13370: out <= 16'h04D6;    16'd13371: out <= 16'h0065;
    16'd13372: out <= 16'h02A8;    16'd13373: out <= 16'h0657;    16'd13374: out <= 16'h0756;    16'd13375: out <= 16'h05D6;
    16'd13376: out <= 16'h0108;    16'd13377: out <= 16'hFFD3;    16'd13378: out <= 16'h0695;    16'd13379: out <= 16'hFE87;
    16'd13380: out <= 16'hFD1A;    16'd13381: out <= 16'hFA18;    16'd13382: out <= 16'h02D5;    16'd13383: out <= 16'h0078;
    16'd13384: out <= 16'h0CC7;    16'd13385: out <= 16'h0083;    16'd13386: out <= 16'h0C08;    16'd13387: out <= 16'h090F;
    16'd13388: out <= 16'hFBB4;    16'd13389: out <= 16'h0437;    16'd13390: out <= 16'h0610;    16'd13391: out <= 16'h0938;
    16'd13392: out <= 16'h0578;    16'd13393: out <= 16'hF8E1;    16'd13394: out <= 16'h09DC;    16'd13395: out <= 16'h083E;
    16'd13396: out <= 16'h02D9;    16'd13397: out <= 16'hFF74;    16'd13398: out <= 16'h00DF;    16'd13399: out <= 16'h027F;
    16'd13400: out <= 16'h0BE6;    16'd13401: out <= 16'hFFD5;    16'd13402: out <= 16'h038A;    16'd13403: out <= 16'h0799;
    16'd13404: out <= 16'h0173;    16'd13405: out <= 16'h01B5;    16'd13406: out <= 16'h0766;    16'd13407: out <= 16'h0409;
    16'd13408: out <= 16'hFCB2;    16'd13409: out <= 16'hFF3E;    16'd13410: out <= 16'h0308;    16'd13411: out <= 16'h0008;
    16'd13412: out <= 16'hFFED;    16'd13413: out <= 16'h005C;    16'd13414: out <= 16'h0726;    16'd13415: out <= 16'h009F;
    16'd13416: out <= 16'h028D;    16'd13417: out <= 16'h008F;    16'd13418: out <= 16'h00D1;    16'd13419: out <= 16'hF7D8;
    16'd13420: out <= 16'hFDB3;    16'd13421: out <= 16'h0475;    16'd13422: out <= 16'h023A;    16'd13423: out <= 16'h04D2;
    16'd13424: out <= 16'h0665;    16'd13425: out <= 16'hFF1A;    16'd13426: out <= 16'h0923;    16'd13427: out <= 16'h02BC;
    16'd13428: out <= 16'h0356;    16'd13429: out <= 16'h029E;    16'd13430: out <= 16'h05A7;    16'd13431: out <= 16'hFF4B;
    16'd13432: out <= 16'h01D8;    16'd13433: out <= 16'h03C3;    16'd13434: out <= 16'h041F;    16'd13435: out <= 16'h0866;
    16'd13436: out <= 16'h0300;    16'd13437: out <= 16'h0283;    16'd13438: out <= 16'h0026;    16'd13439: out <= 16'h03AB;
    16'd13440: out <= 16'h0B7B;    16'd13441: out <= 16'hFDD1;    16'd13442: out <= 16'h0690;    16'd13443: out <= 16'h04B9;
    16'd13444: out <= 16'h0166;    16'd13445: out <= 16'h01C8;    16'd13446: out <= 16'h0231;    16'd13447: out <= 16'h091A;
    16'd13448: out <= 16'h0334;    16'd13449: out <= 16'h066F;    16'd13450: out <= 16'h0377;    16'd13451: out <= 16'h0432;
    16'd13452: out <= 16'h01DC;    16'd13453: out <= 16'h0271;    16'd13454: out <= 16'h0455;    16'd13455: out <= 16'h04BB;
    16'd13456: out <= 16'hFF48;    16'd13457: out <= 16'h0654;    16'd13458: out <= 16'h00FE;    16'd13459: out <= 16'h00D3;
    16'd13460: out <= 16'h0456;    16'd13461: out <= 16'h09AF;    16'd13462: out <= 16'h011B;    16'd13463: out <= 16'hFEC1;
    16'd13464: out <= 16'h0452;    16'd13465: out <= 16'h0744;    16'd13466: out <= 16'h08C6;    16'd13467: out <= 16'h0618;
    16'd13468: out <= 16'h036C;    16'd13469: out <= 16'h0276;    16'd13470: out <= 16'hFC27;    16'd13471: out <= 16'hFC88;
    16'd13472: out <= 16'h0364;    16'd13473: out <= 16'h029C;    16'd13474: out <= 16'h0000;    16'd13475: out <= 16'hFC59;
    16'd13476: out <= 16'h063F;    16'd13477: out <= 16'hFFB8;    16'd13478: out <= 16'h029A;    16'd13479: out <= 16'h028D;
    16'd13480: out <= 16'h051D;    16'd13481: out <= 16'h0999;    16'd13482: out <= 16'h062D;    16'd13483: out <= 16'h0642;
    16'd13484: out <= 16'h05CB;    16'd13485: out <= 16'h0650;    16'd13486: out <= 16'h098E;    16'd13487: out <= 16'h0B12;
    16'd13488: out <= 16'h0295;    16'd13489: out <= 16'h0415;    16'd13490: out <= 16'hFF61;    16'd13491: out <= 16'h00CA;
    16'd13492: out <= 16'h01E3;    16'd13493: out <= 16'h0128;    16'd13494: out <= 16'h0310;    16'd13495: out <= 16'hFFF8;
    16'd13496: out <= 16'h002B;    16'd13497: out <= 16'hFEA5;    16'd13498: out <= 16'h0A7E;    16'd13499: out <= 16'h0205;
    16'd13500: out <= 16'h05B2;    16'd13501: out <= 16'h0592;    16'd13502: out <= 16'h0274;    16'd13503: out <= 16'h005B;
    16'd13504: out <= 16'h00A2;    16'd13505: out <= 16'h0516;    16'd13506: out <= 16'h05C1;    16'd13507: out <= 16'hFE4A;
    16'd13508: out <= 16'h0504;    16'd13509: out <= 16'h02AD;    16'd13510: out <= 16'h06CA;    16'd13511: out <= 16'h0261;
    16'd13512: out <= 16'h0545;    16'd13513: out <= 16'h0903;    16'd13514: out <= 16'h0382;    16'd13515: out <= 16'h03B5;
    16'd13516: out <= 16'h05B8;    16'd13517: out <= 16'h02ED;    16'd13518: out <= 16'h0776;    16'd13519: out <= 16'hFD1E;
    16'd13520: out <= 16'h0000;    16'd13521: out <= 16'h0B1E;    16'd13522: out <= 16'h0329;    16'd13523: out <= 16'h06F1;
    16'd13524: out <= 16'h05B3;    16'd13525: out <= 16'h000E;    16'd13526: out <= 16'h024F;    16'd13527: out <= 16'h06D4;
    16'd13528: out <= 16'h00DF;    16'd13529: out <= 16'h0482;    16'd13530: out <= 16'hFE5F;    16'd13531: out <= 16'hFFEF;
    16'd13532: out <= 16'h01E1;    16'd13533: out <= 16'hFB29;    16'd13534: out <= 16'hFEB3;    16'd13535: out <= 16'h021E;
    16'd13536: out <= 16'hFDA7;    16'd13537: out <= 16'hFE88;    16'd13538: out <= 16'h014F;    16'd13539: out <= 16'h024B;
    16'd13540: out <= 16'hFCEB;    16'd13541: out <= 16'hFFC5;    16'd13542: out <= 16'hFBB8;    16'd13543: out <= 16'hFAD8;
    16'd13544: out <= 16'hFC6A;    16'd13545: out <= 16'h0062;    16'd13546: out <= 16'h01D4;    16'd13547: out <= 16'h0149;
    16'd13548: out <= 16'hFF31;    16'd13549: out <= 16'h006C;    16'd13550: out <= 16'hFC87;    16'd13551: out <= 16'h02B2;
    16'd13552: out <= 16'hFE3B;    16'd13553: out <= 16'hFFCA;    16'd13554: out <= 16'h034F;    16'd13555: out <= 16'h021B;
    16'd13556: out <= 16'h0446;    16'd13557: out <= 16'hF97B;    16'd13558: out <= 16'hFBCB;    16'd13559: out <= 16'hF7F8;
    16'd13560: out <= 16'hFD65;    16'd13561: out <= 16'hFCC2;    16'd13562: out <= 16'hFFF5;    16'd13563: out <= 16'hF8A7;
    16'd13564: out <= 16'hFF51;    16'd13565: out <= 16'hFC4A;    16'd13566: out <= 16'h01F9;    16'd13567: out <= 16'h034C;
    16'd13568: out <= 16'hFAF8;    16'd13569: out <= 16'hFEB3;    16'd13570: out <= 16'h0181;    16'd13571: out <= 16'hFF17;
    16'd13572: out <= 16'h007C;    16'd13573: out <= 16'hFAEF;    16'd13574: out <= 16'h04F9;    16'd13575: out <= 16'h00CB;
    16'd13576: out <= 16'h034F;    16'd13577: out <= 16'hFE9F;    16'd13578: out <= 16'h02A7;    16'd13579: out <= 16'hFF12;
    16'd13580: out <= 16'hFADC;    16'd13581: out <= 16'h044E;    16'd13582: out <= 16'h036C;    16'd13583: out <= 16'hF738;
    16'd13584: out <= 16'hF7FB;    16'd13585: out <= 16'h018D;    16'd13586: out <= 16'hFC59;    16'd13587: out <= 16'hFA17;
    16'd13588: out <= 16'h00B8;    16'd13589: out <= 16'hFB06;    16'd13590: out <= 16'hFB0F;    16'd13591: out <= 16'h00CA;
    16'd13592: out <= 16'hFD3B;    16'd13593: out <= 16'h0505;    16'd13594: out <= 16'h0653;    16'd13595: out <= 16'h0673;
    16'd13596: out <= 16'h0A10;    16'd13597: out <= 16'h018F;    16'd13598: out <= 16'hFCDE;    16'd13599: out <= 16'hFBB3;
    16'd13600: out <= 16'hFF38;    16'd13601: out <= 16'h0017;    16'd13602: out <= 16'h09A8;    16'd13603: out <= 16'h04E7;
    16'd13604: out <= 16'h05D8;    16'd13605: out <= 16'h02E8;    16'd13606: out <= 16'h064F;    16'd13607: out <= 16'hFD65;
    16'd13608: out <= 16'h013F;    16'd13609: out <= 16'h02C6;    16'd13610: out <= 16'h08BD;    16'd13611: out <= 16'h071D;
    16'd13612: out <= 16'h0AA8;    16'd13613: out <= 16'h03C7;    16'd13614: out <= 16'h042A;    16'd13615: out <= 16'h0431;
    16'd13616: out <= 16'hFE68;    16'd13617: out <= 16'h032D;    16'd13618: out <= 16'h003A;    16'd13619: out <= 16'h019C;
    16'd13620: out <= 16'h0036;    16'd13621: out <= 16'h0056;    16'd13622: out <= 16'h05C5;    16'd13623: out <= 16'h04E2;
    16'd13624: out <= 16'h0806;    16'd13625: out <= 16'h04F7;    16'd13626: out <= 16'h00DE;    16'd13627: out <= 16'h0926;
    16'd13628: out <= 16'h06B8;    16'd13629: out <= 16'h08EC;    16'd13630: out <= 16'h00FC;    16'd13631: out <= 16'hFE90;
    16'd13632: out <= 16'h0A17;    16'd13633: out <= 16'h0BBE;    16'd13634: out <= 16'h03ED;    16'd13635: out <= 16'hFF8B;
    16'd13636: out <= 16'h01E9;    16'd13637: out <= 16'h052E;    16'd13638: out <= 16'h0402;    16'd13639: out <= 16'h0176;
    16'd13640: out <= 16'h03CE;    16'd13641: out <= 16'h0403;    16'd13642: out <= 16'h07B7;    16'd13643: out <= 16'h05E4;
    16'd13644: out <= 16'h04E7;    16'd13645: out <= 16'h0625;    16'd13646: out <= 16'h081B;    16'd13647: out <= 16'hFCED;
    16'd13648: out <= 16'h005F;    16'd13649: out <= 16'h01D3;    16'd13650: out <= 16'h0318;    16'd13651: out <= 16'h047B;
    16'd13652: out <= 16'h03AB;    16'd13653: out <= 16'h005E;    16'd13654: out <= 16'h07B4;    16'd13655: out <= 16'h04AE;
    16'd13656: out <= 16'h0352;    16'd13657: out <= 16'h033E;    16'd13658: out <= 16'h0695;    16'd13659: out <= 16'hFB8A;
    16'd13660: out <= 16'h0174;    16'd13661: out <= 16'h0152;    16'd13662: out <= 16'h0619;    16'd13663: out <= 16'hFF41;
    16'd13664: out <= 16'h0003;    16'd13665: out <= 16'h06D1;    16'd13666: out <= 16'h013C;    16'd13667: out <= 16'hFD1F;
    16'd13668: out <= 16'h01A9;    16'd13669: out <= 16'hFF4C;    16'd13670: out <= 16'h002B;    16'd13671: out <= 16'h087A;
    16'd13672: out <= 16'h0387;    16'd13673: out <= 16'h04BC;    16'd13674: out <= 16'h070F;    16'd13675: out <= 16'h00B6;
    16'd13676: out <= 16'h023E;    16'd13677: out <= 16'h0624;    16'd13678: out <= 16'hFF16;    16'd13679: out <= 16'h0010;
    16'd13680: out <= 16'h04E5;    16'd13681: out <= 16'h04C7;    16'd13682: out <= 16'hFF4E;    16'd13683: out <= 16'h0D41;
    16'd13684: out <= 16'h0212;    16'd13685: out <= 16'h0680;    16'd13686: out <= 16'h0532;    16'd13687: out <= 16'h0098;
    16'd13688: out <= 16'h0210;    16'd13689: out <= 16'h03C0;    16'd13690: out <= 16'hFD96;    16'd13691: out <= 16'h0376;
    16'd13692: out <= 16'h0249;    16'd13693: out <= 16'h031A;    16'd13694: out <= 16'h04F8;    16'd13695: out <= 16'hFF3C;
    16'd13696: out <= 16'h0099;    16'd13697: out <= 16'h046A;    16'd13698: out <= 16'h0BDD;    16'd13699: out <= 16'h0474;
    16'd13700: out <= 16'h0940;    16'd13701: out <= 16'h09DC;    16'd13702: out <= 16'h06EA;    16'd13703: out <= 16'h00F2;
    16'd13704: out <= 16'h0317;    16'd13705: out <= 16'h08C1;    16'd13706: out <= 16'h04E4;    16'd13707: out <= 16'h049C;
    16'd13708: out <= 16'h0333;    16'd13709: out <= 16'h00C8;    16'd13710: out <= 16'h0207;    16'd13711: out <= 16'hFFDC;
    16'd13712: out <= 16'h00A3;    16'd13713: out <= 16'h04B2;    16'd13714: out <= 16'h0AFD;    16'd13715: out <= 16'h0444;
    16'd13716: out <= 16'h015E;    16'd13717: out <= 16'h0628;    16'd13718: out <= 16'h001C;    16'd13719: out <= 16'h01D9;
    16'd13720: out <= 16'h0157;    16'd13721: out <= 16'h10A6;    16'd13722: out <= 16'h074B;    16'd13723: out <= 16'hFBA9;
    16'd13724: out <= 16'h05DB;    16'd13725: out <= 16'h050D;    16'd13726: out <= 16'h03C8;    16'd13727: out <= 16'h038C;
    16'd13728: out <= 16'h0370;    16'd13729: out <= 16'h0CB2;    16'd13730: out <= 16'hFB9A;    16'd13731: out <= 16'h00FF;
    16'd13732: out <= 16'h0848;    16'd13733: out <= 16'h0956;    16'd13734: out <= 16'h0439;    16'd13735: out <= 16'h0880;
    16'd13736: out <= 16'hFE02;    16'd13737: out <= 16'h035A;    16'd13738: out <= 16'h062B;    16'd13739: out <= 16'h01B6;
    16'd13740: out <= 16'h01F5;    16'd13741: out <= 16'h021B;    16'd13742: out <= 16'h057C;    16'd13743: out <= 16'h02CA;
    16'd13744: out <= 16'h022A;    16'd13745: out <= 16'h0212;    16'd13746: out <= 16'h042B;    16'd13747: out <= 16'h05CB;
    16'd13748: out <= 16'h0101;    16'd13749: out <= 16'hFC32;    16'd13750: out <= 16'hFDFE;    16'd13751: out <= 16'hFE3C;
    16'd13752: out <= 16'h078D;    16'd13753: out <= 16'h092C;    16'd13754: out <= 16'h050C;    16'd13755: out <= 16'h0386;
    16'd13756: out <= 16'h021D;    16'd13757: out <= 16'h002A;    16'd13758: out <= 16'hFE7C;    16'd13759: out <= 16'h0122;
    16'd13760: out <= 16'h009C;    16'd13761: out <= 16'hFEBB;    16'd13762: out <= 16'h026B;    16'd13763: out <= 16'h0EA4;
    16'd13764: out <= 16'h0632;    16'd13765: out <= 16'h0656;    16'd13766: out <= 16'h008E;    16'd13767: out <= 16'hFC06;
    16'd13768: out <= 16'h0370;    16'd13769: out <= 16'h066D;    16'd13770: out <= 16'h057D;    16'd13771: out <= 16'h0610;
    16'd13772: out <= 16'h0613;    16'd13773: out <= 16'hFE6E;    16'd13774: out <= 16'h054B;    16'd13775: out <= 16'h063C;
    16'd13776: out <= 16'hFEEB;    16'd13777: out <= 16'h0411;    16'd13778: out <= 16'h04FD;    16'd13779: out <= 16'h04BB;
    16'd13780: out <= 16'h0590;    16'd13781: out <= 16'h00F4;    16'd13782: out <= 16'hFBE2;    16'd13783: out <= 16'hFDDE;
    16'd13784: out <= 16'hFFB8;    16'd13785: out <= 16'hFEF4;    16'd13786: out <= 16'h04E1;    16'd13787: out <= 16'h01B5;
    16'd13788: out <= 16'hFFBF;    16'd13789: out <= 16'hFB60;    16'd13790: out <= 16'hF9EE;    16'd13791: out <= 16'hFF5B;
    16'd13792: out <= 16'h00DC;    16'd13793: out <= 16'hFCC2;    16'd13794: out <= 16'hFB7F;    16'd13795: out <= 16'h04A0;
    16'd13796: out <= 16'hFBA9;    16'd13797: out <= 16'h04F0;    16'd13798: out <= 16'hFD3B;    16'd13799: out <= 16'hFC64;
    16'd13800: out <= 16'h00DA;    16'd13801: out <= 16'h046E;    16'd13802: out <= 16'hFA0D;    16'd13803: out <= 16'hFC36;
    16'd13804: out <= 16'h0180;    16'd13805: out <= 16'h049E;    16'd13806: out <= 16'hFF5E;    16'd13807: out <= 16'hFF50;
    16'd13808: out <= 16'hFCD8;    16'd13809: out <= 16'h00C7;    16'd13810: out <= 16'hFCBE;    16'd13811: out <= 16'h0181;
    16'd13812: out <= 16'hFA65;    16'd13813: out <= 16'h059A;    16'd13814: out <= 16'h0394;    16'd13815: out <= 16'h0234;
    16'd13816: out <= 16'hFCFF;    16'd13817: out <= 16'h020B;    16'd13818: out <= 16'h020B;    16'd13819: out <= 16'hFE90;
    16'd13820: out <= 16'hFD38;    16'd13821: out <= 16'hFD0A;    16'd13822: out <= 16'h0361;    16'd13823: out <= 16'hF9FB;
    16'd13824: out <= 16'hF6BA;    16'd13825: out <= 16'h0138;    16'd13826: out <= 16'hF641;    16'd13827: out <= 16'hFF28;
    16'd13828: out <= 16'h0434;    16'd13829: out <= 16'hFE18;    16'd13830: out <= 16'h036C;    16'd13831: out <= 16'h007F;
    16'd13832: out <= 16'hF4B9;    16'd13833: out <= 16'hFD20;    16'd13834: out <= 16'hFF02;    16'd13835: out <= 16'hFF7E;
    16'd13836: out <= 16'hFF81;    16'd13837: out <= 16'hF751;    16'd13838: out <= 16'h089A;    16'd13839: out <= 16'h02A6;
    16'd13840: out <= 16'h057C;    16'd13841: out <= 16'hFD34;    16'd13842: out <= 16'hFFA5;    16'd13843: out <= 16'hFAE5;
    16'd13844: out <= 16'hFE9D;    16'd13845: out <= 16'h0591;    16'd13846: out <= 16'hFC4B;    16'd13847: out <= 16'h0125;
    16'd13848: out <= 16'h0359;    16'd13849: out <= 16'hFDE1;    16'd13850: out <= 16'hFD2C;    16'd13851: out <= 16'hFB91;
    16'd13852: out <= 16'hFED0;    16'd13853: out <= 16'h035C;    16'd13854: out <= 16'h0319;    16'd13855: out <= 16'hFC1F;
    16'd13856: out <= 16'hFEA6;    16'd13857: out <= 16'h087D;    16'd13858: out <= 16'h035E;    16'd13859: out <= 16'h0164;
    16'd13860: out <= 16'h0325;    16'd13861: out <= 16'h0948;    16'd13862: out <= 16'hFF0C;    16'd13863: out <= 16'h0354;
    16'd13864: out <= 16'h010F;    16'd13865: out <= 16'h03BF;    16'd13866: out <= 16'h01EC;    16'd13867: out <= 16'h05BE;
    16'd13868: out <= 16'h06AF;    16'd13869: out <= 16'h02D3;    16'd13870: out <= 16'h047F;    16'd13871: out <= 16'h02BF;
    16'd13872: out <= 16'h091B;    16'd13873: out <= 16'h03FF;    16'd13874: out <= 16'h0B0E;    16'd13875: out <= 16'h038C;
    16'd13876: out <= 16'h0474;    16'd13877: out <= 16'h00A0;    16'd13878: out <= 16'h079C;    16'd13879: out <= 16'h0A35;
    16'd13880: out <= 16'h0745;    16'd13881: out <= 16'hFE05;    16'd13882: out <= 16'h004B;    16'd13883: out <= 16'hFB6A;
    16'd13884: out <= 16'h0055;    16'd13885: out <= 16'h06B7;    16'd13886: out <= 16'h0018;    16'd13887: out <= 16'h00E1;
    16'd13888: out <= 16'h091D;    16'd13889: out <= 16'h065A;    16'd13890: out <= 16'h0134;    16'd13891: out <= 16'h019C;
    16'd13892: out <= 16'h02A5;    16'd13893: out <= 16'h0791;    16'd13894: out <= 16'hFC92;    16'd13895: out <= 16'hFF09;
    16'd13896: out <= 16'hFDF4;    16'd13897: out <= 16'h0E7E;    16'd13898: out <= 16'h01D9;    16'd13899: out <= 16'h05F4;
    16'd13900: out <= 16'h0680;    16'd13901: out <= 16'h02D0;    16'd13902: out <= 16'h038E;    16'd13903: out <= 16'h0360;
    16'd13904: out <= 16'hFF1F;    16'd13905: out <= 16'h02D5;    16'd13906: out <= 16'h06FE;    16'd13907: out <= 16'h00B8;
    16'd13908: out <= 16'h06E1;    16'd13909: out <= 16'hFE7F;    16'd13910: out <= 16'h0875;    16'd13911: out <= 16'h01B8;
    16'd13912: out <= 16'h01FC;    16'd13913: out <= 16'h0664;    16'd13914: out <= 16'hF8FC;    16'd13915: out <= 16'h0983;
    16'd13916: out <= 16'h02E0;    16'd13917: out <= 16'h056E;    16'd13918: out <= 16'hFE0C;    16'd13919: out <= 16'h050E;
    16'd13920: out <= 16'h02AF;    16'd13921: out <= 16'h0533;    16'd13922: out <= 16'h0818;    16'd13923: out <= 16'h04C2;
    16'd13924: out <= 16'h01AC;    16'd13925: out <= 16'h024E;    16'd13926: out <= 16'h0204;    16'd13927: out <= 16'h0228;
    16'd13928: out <= 16'h0341;    16'd13929: out <= 16'h0746;    16'd13930: out <= 16'h0262;    16'd13931: out <= 16'hFDD1;
    16'd13932: out <= 16'h0398;    16'd13933: out <= 16'h053E;    16'd13934: out <= 16'h08D2;    16'd13935: out <= 16'h0809;
    16'd13936: out <= 16'h05AB;    16'd13937: out <= 16'h009F;    16'd13938: out <= 16'h0425;    16'd13939: out <= 16'h00A9;
    16'd13940: out <= 16'h04AE;    16'd13941: out <= 16'h020A;    16'd13942: out <= 16'hFE9D;    16'd13943: out <= 16'hFE4D;
    16'd13944: out <= 16'h0A22;    16'd13945: out <= 16'h0309;    16'd13946: out <= 16'h0A42;    16'd13947: out <= 16'h072F;
    16'd13948: out <= 16'h04BB;    16'd13949: out <= 16'hFF36;    16'd13950: out <= 16'h0085;    16'd13951: out <= 16'h0482;
    16'd13952: out <= 16'h01EA;    16'd13953: out <= 16'h003D;    16'd13954: out <= 16'h05FA;    16'd13955: out <= 16'h0B85;
    16'd13956: out <= 16'h09AB;    16'd13957: out <= 16'hFC68;    16'd13958: out <= 16'h0812;    16'd13959: out <= 16'h08CA;
    16'd13960: out <= 16'h0362;    16'd13961: out <= 16'hFED1;    16'd13962: out <= 16'h0416;    16'd13963: out <= 16'h06C9;
    16'd13964: out <= 16'h0873;    16'd13965: out <= 16'h0098;    16'd13966: out <= 16'h00D5;    16'd13967: out <= 16'h07CE;
    16'd13968: out <= 16'h01FD;    16'd13969: out <= 16'h0543;    16'd13970: out <= 16'h027D;    16'd13971: out <= 16'hFFE1;
    16'd13972: out <= 16'h0AD7;    16'd13973: out <= 16'h0064;    16'd13974: out <= 16'h017A;    16'd13975: out <= 16'hFB7A;
    16'd13976: out <= 16'h04D0;    16'd13977: out <= 16'hFC3F;    16'd13978: out <= 16'hFD5D;    16'd13979: out <= 16'h010B;
    16'd13980: out <= 16'h042C;    16'd13981: out <= 16'h066B;    16'd13982: out <= 16'h03F7;    16'd13983: out <= 16'h04FF;
    16'd13984: out <= 16'h0712;    16'd13985: out <= 16'h018F;    16'd13986: out <= 16'h024D;    16'd13987: out <= 16'h039D;
    16'd13988: out <= 16'h06B5;    16'd13989: out <= 16'h0112;    16'd13990: out <= 16'h030E;    16'd13991: out <= 16'h0393;
    16'd13992: out <= 16'h06A5;    16'd13993: out <= 16'h0219;    16'd13994: out <= 16'h0A84;    16'd13995: out <= 16'h0DB3;
    16'd13996: out <= 16'h084E;    16'd13997: out <= 16'h04FA;    16'd13998: out <= 16'h089F;    16'd13999: out <= 16'h076A;
    16'd14000: out <= 16'h0380;    16'd14001: out <= 16'hF9F3;    16'd14002: out <= 16'h01A6;    16'd14003: out <= 16'hFE23;
    16'd14004: out <= 16'h0312;    16'd14005: out <= 16'h07AB;    16'd14006: out <= 16'h02C0;    16'd14007: out <= 16'h01BC;
    16'd14008: out <= 16'h0227;    16'd14009: out <= 16'h0353;    16'd14010: out <= 16'h01F0;    16'd14011: out <= 16'h0170;
    16'd14012: out <= 16'h054D;    16'd14013: out <= 16'hFE07;    16'd14014: out <= 16'h052C;    16'd14015: out <= 16'h00F1;
    16'd14016: out <= 16'hFD26;    16'd14017: out <= 16'h0617;    16'd14018: out <= 16'h0473;    16'd14019: out <= 16'h0707;
    16'd14020: out <= 16'h0428;    16'd14021: out <= 16'h041C;    16'd14022: out <= 16'h05DE;    16'd14023: out <= 16'h012A;
    16'd14024: out <= 16'h076E;    16'd14025: out <= 16'hFB90;    16'd14026: out <= 16'h00C5;    16'd14027: out <= 16'hFCA7;
    16'd14028: out <= 16'h05B2;    16'd14029: out <= 16'h02C9;    16'd14030: out <= 16'h0459;    16'd14031: out <= 16'h0600;
    16'd14032: out <= 16'h03FE;    16'd14033: out <= 16'h076A;    16'd14034: out <= 16'h0126;    16'd14035: out <= 16'h061A;
    16'd14036: out <= 16'hFEE1;    16'd14037: out <= 16'h00EC;    16'd14038: out <= 16'h003B;    16'd14039: out <= 16'hFEEF;
    16'd14040: out <= 16'h042A;    16'd14041: out <= 16'hFA3D;    16'd14042: out <= 16'hFFEF;    16'd14043: out <= 16'h0074;
    16'd14044: out <= 16'h0307;    16'd14045: out <= 16'h0076;    16'd14046: out <= 16'h0131;    16'd14047: out <= 16'hFD09;
    16'd14048: out <= 16'h0402;    16'd14049: out <= 16'h00BC;    16'd14050: out <= 16'h0088;    16'd14051: out <= 16'hFCA8;
    16'd14052: out <= 16'h023D;    16'd14053: out <= 16'hFA8B;    16'd14054: out <= 16'hFF56;    16'd14055: out <= 16'h010E;
    16'd14056: out <= 16'hFFCD;    16'd14057: out <= 16'hF771;    16'd14058: out <= 16'hFC34;    16'd14059: out <= 16'h012C;
    16'd14060: out <= 16'hFE2D;    16'd14061: out <= 16'hF9DB;    16'd14062: out <= 16'h077D;    16'd14063: out <= 16'hFFF1;
    16'd14064: out <= 16'h0071;    16'd14065: out <= 16'h0154;    16'd14066: out <= 16'hFED9;    16'd14067: out <= 16'h0339;
    16'd14068: out <= 16'hFFE6;    16'd14069: out <= 16'hFE52;    16'd14070: out <= 16'hF619;    16'd14071: out <= 16'h01DC;
    16'd14072: out <= 16'h04BB;    16'd14073: out <= 16'h0200;    16'd14074: out <= 16'h00DB;    16'd14075: out <= 16'hFCAF;
    16'd14076: out <= 16'hFF05;    16'd14077: out <= 16'h0199;    16'd14078: out <= 16'h003F;    16'd14079: out <= 16'hF830;
    16'd14080: out <= 16'hFDCE;    16'd14081: out <= 16'h043C;    16'd14082: out <= 16'h023A;    16'd14083: out <= 16'hFF33;
    16'd14084: out <= 16'h03B6;    16'd14085: out <= 16'hFA03;    16'd14086: out <= 16'hFE6C;    16'd14087: out <= 16'hF98F;
    16'd14088: out <= 16'h042B;    16'd14089: out <= 16'h0097;    16'd14090: out <= 16'hFF63;    16'd14091: out <= 16'hFF8C;
    16'd14092: out <= 16'h0314;    16'd14093: out <= 16'hFED9;    16'd14094: out <= 16'hFBFD;    16'd14095: out <= 16'h034D;
    16'd14096: out <= 16'hFCE6;    16'd14097: out <= 16'h068C;    16'd14098: out <= 16'hF9A2;    16'd14099: out <= 16'hFEDD;
    16'd14100: out <= 16'h004D;    16'd14101: out <= 16'h032A;    16'd14102: out <= 16'h0724;    16'd14103: out <= 16'hFE44;
    16'd14104: out <= 16'hF5E9;    16'd14105: out <= 16'h01D4;    16'd14106: out <= 16'h0063;    16'd14107: out <= 16'hFC40;
    16'd14108: out <= 16'h04C3;    16'd14109: out <= 16'hFE4B;    16'd14110: out <= 16'hFF7B;    16'd14111: out <= 16'h0A08;
    16'd14112: out <= 16'hFBDD;    16'd14113: out <= 16'hFDD2;    16'd14114: out <= 16'h0411;    16'd14115: out <= 16'h041B;
    16'd14116: out <= 16'hFCFC;    16'd14117: out <= 16'h069B;    16'd14118: out <= 16'h053A;    16'd14119: out <= 16'h0036;
    16'd14120: out <= 16'h05AD;    16'd14121: out <= 16'h0306;    16'd14122: out <= 16'h03A7;    16'd14123: out <= 16'h0A98;
    16'd14124: out <= 16'h058C;    16'd14125: out <= 16'h0CBA;    16'd14126: out <= 16'h06EB;    16'd14127: out <= 16'hFD16;
    16'd14128: out <= 16'h0919;    16'd14129: out <= 16'h045D;    16'd14130: out <= 16'h00F9;    16'd14131: out <= 16'h0476;
    16'd14132: out <= 16'h04F1;    16'd14133: out <= 16'h0560;    16'd14134: out <= 16'h07B2;    16'd14135: out <= 16'h0399;
    16'd14136: out <= 16'h009B;    16'd14137: out <= 16'h01A3;    16'd14138: out <= 16'h0635;    16'd14139: out <= 16'hFFAF;
    16'd14140: out <= 16'h0484;    16'd14141: out <= 16'h0D38;    16'd14142: out <= 16'h026A;    16'd14143: out <= 16'h07A5;
    16'd14144: out <= 16'h04A8;    16'd14145: out <= 16'h0715;    16'd14146: out <= 16'h0502;    16'd14147: out <= 16'h04B0;
    16'd14148: out <= 16'hFF29;    16'd14149: out <= 16'h0041;    16'd14150: out <= 16'h06A5;    16'd14151: out <= 16'h06DB;
    16'd14152: out <= 16'h0832;    16'd14153: out <= 16'h0808;    16'd14154: out <= 16'h0299;    16'd14155: out <= 16'h0416;
    16'd14156: out <= 16'hFFC0;    16'd14157: out <= 16'h00F2;    16'd14158: out <= 16'h0302;    16'd14159: out <= 16'h0199;
    16'd14160: out <= 16'h05FD;    16'd14161: out <= 16'h0AC0;    16'd14162: out <= 16'h0386;    16'd14163: out <= 16'h0031;
    16'd14164: out <= 16'h0441;    16'd14165: out <= 16'hFEE1;    16'd14166: out <= 16'h0424;    16'd14167: out <= 16'h0085;
    16'd14168: out <= 16'h0109;    16'd14169: out <= 16'hFE6F;    16'd14170: out <= 16'h0052;    16'd14171: out <= 16'h0183;
    16'd14172: out <= 16'h05B7;    16'd14173: out <= 16'hFDDD;    16'd14174: out <= 16'h0417;    16'd14175: out <= 16'h060C;
    16'd14176: out <= 16'h0E6B;    16'd14177: out <= 16'hFEFC;    16'd14178: out <= 16'h0088;    16'd14179: out <= 16'h020F;
    16'd14180: out <= 16'h0274;    16'd14181: out <= 16'h05D6;    16'd14182: out <= 16'h02C5;    16'd14183: out <= 16'h0454;
    16'd14184: out <= 16'h028B;    16'd14185: out <= 16'h02A9;    16'd14186: out <= 16'h07BE;    16'd14187: out <= 16'h01FA;
    16'd14188: out <= 16'h01E1;    16'd14189: out <= 16'h0CD1;    16'd14190: out <= 16'h09CE;    16'd14191: out <= 16'h0A86;
    16'd14192: out <= 16'h0225;    16'd14193: out <= 16'h0325;    16'd14194: out <= 16'h052C;    16'd14195: out <= 16'h07DD;
    16'd14196: out <= 16'h0214;    16'd14197: out <= 16'h0E16;    16'd14198: out <= 16'h0350;    16'd14199: out <= 16'hFE33;
    16'd14200: out <= 16'h0283;    16'd14201: out <= 16'h02C8;    16'd14202: out <= 16'h041F;    16'd14203: out <= 16'hFF26;
    16'd14204: out <= 16'h0271;    16'd14205: out <= 16'h0BFB;    16'd14206: out <= 16'h049B;    16'd14207: out <= 16'h07E4;
    16'd14208: out <= 16'h03C7;    16'd14209: out <= 16'h03E7;    16'd14210: out <= 16'h041A;    16'd14211: out <= 16'h0455;
    16'd14212: out <= 16'hFFC8;    16'd14213: out <= 16'h06FF;    16'd14214: out <= 16'hFCA3;    16'd14215: out <= 16'hFE71;
    16'd14216: out <= 16'h080E;    16'd14217: out <= 16'h0333;    16'd14218: out <= 16'h0805;    16'd14219: out <= 16'hFE4F;
    16'd14220: out <= 16'h08CD;    16'd14221: out <= 16'hFE36;    16'd14222: out <= 16'h01E0;    16'd14223: out <= 16'h0313;
    16'd14224: out <= 16'hFCE7;    16'd14225: out <= 16'h0782;    16'd14226: out <= 16'h0307;    16'd14227: out <= 16'h09C6;
    16'd14228: out <= 16'h0246;    16'd14229: out <= 16'h0247;    16'd14230: out <= 16'hF9E8;    16'd14231: out <= 16'h02C1;
    16'd14232: out <= 16'h03FC;    16'd14233: out <= 16'hFF7A;    16'd14234: out <= 16'h0603;    16'd14235: out <= 16'h05D2;
    16'd14236: out <= 16'h0090;    16'd14237: out <= 16'hFF2B;    16'd14238: out <= 16'hFAE6;    16'd14239: out <= 16'h064A;
    16'd14240: out <= 16'h010A;    16'd14241: out <= 16'h063A;    16'd14242: out <= 16'h0589;    16'd14243: out <= 16'h0A37;
    16'd14244: out <= 16'h05AB;    16'd14245: out <= 16'hFFC5;    16'd14246: out <= 16'h001F;    16'd14247: out <= 16'h0441;
    16'd14248: out <= 16'h014E;    16'd14249: out <= 16'h00CB;    16'd14250: out <= 16'h051A;    16'd14251: out <= 16'hFF68;
    16'd14252: out <= 16'h099A;    16'd14253: out <= 16'hF9DF;    16'd14254: out <= 16'h0733;    16'd14255: out <= 16'h01A1;
    16'd14256: out <= 16'h02EB;    16'd14257: out <= 16'h0AAE;    16'd14258: out <= 16'h00AD;    16'd14259: out <= 16'h0421;
    16'd14260: out <= 16'hFE53;    16'd14261: out <= 16'h031B;    16'd14262: out <= 16'h053D;    16'd14263: out <= 16'h0345;
    16'd14264: out <= 16'h0452;    16'd14265: out <= 16'h06EE;    16'd14266: out <= 16'hFBF1;    16'd14267: out <= 16'h0601;
    16'd14268: out <= 16'h0579;    16'd14269: out <= 16'h0196;    16'd14270: out <= 16'h07AC;    16'd14271: out <= 16'h0372;
    16'd14272: out <= 16'h047B;    16'd14273: out <= 16'h0298;    16'd14274: out <= 16'hFC42;    16'd14275: out <= 16'h09E7;
    16'd14276: out <= 16'hFFCA;    16'd14277: out <= 16'h02D4;    16'd14278: out <= 16'h0610;    16'd14279: out <= 16'h01B2;
    16'd14280: out <= 16'h01C1;    16'd14281: out <= 16'h05E8;    16'd14282: out <= 16'h0645;    16'd14283: out <= 16'h0446;
    16'd14284: out <= 16'h0963;    16'd14285: out <= 16'hFFC3;    16'd14286: out <= 16'h0534;    16'd14287: out <= 16'h0052;
    16'd14288: out <= 16'hFFC5;    16'd14289: out <= 16'hFFE6;    16'd14290: out <= 16'hFBB7;    16'd14291: out <= 16'hF7DD;
    16'd14292: out <= 16'hFF3E;    16'd14293: out <= 16'h0986;    16'd14294: out <= 16'h02FD;    16'd14295: out <= 16'h0112;
    16'd14296: out <= 16'h0549;    16'd14297: out <= 16'h084B;    16'd14298: out <= 16'hFC80;    16'd14299: out <= 16'hFF8B;
    16'd14300: out <= 16'h01B0;    16'd14301: out <= 16'h03C5;    16'd14302: out <= 16'h0235;    16'd14303: out <= 16'h0222;
    16'd14304: out <= 16'h0378;    16'd14305: out <= 16'h0045;    16'd14306: out <= 16'hFB08;    16'd14307: out <= 16'h0587;
    16'd14308: out <= 16'hFAD6;    16'd14309: out <= 16'h0407;    16'd14310: out <= 16'h0057;    16'd14311: out <= 16'h0583;
    16'd14312: out <= 16'h07AB;    16'd14313: out <= 16'hF960;    16'd14314: out <= 16'h0360;    16'd14315: out <= 16'hFF91;
    16'd14316: out <= 16'h00CB;    16'd14317: out <= 16'h0768;    16'd14318: out <= 16'hFCB0;    16'd14319: out <= 16'h04EE;
    16'd14320: out <= 16'h00EA;    16'd14321: out <= 16'hFDCB;    16'd14322: out <= 16'hF9E3;    16'd14323: out <= 16'h00A7;
    16'd14324: out <= 16'h00EC;    16'd14325: out <= 16'h01A3;    16'd14326: out <= 16'hFFEA;    16'd14327: out <= 16'hF8A1;
    16'd14328: out <= 16'hFE2A;    16'd14329: out <= 16'hFF9F;    16'd14330: out <= 16'hFFCF;    16'd14331: out <= 16'hFF2A;
    16'd14332: out <= 16'hFD9F;    16'd14333: out <= 16'h0553;    16'd14334: out <= 16'h000C;    16'd14335: out <= 16'h0550;
    16'd14336: out <= 16'h0272;    16'd14337: out <= 16'hFB56;    16'd14338: out <= 16'hFBB0;    16'd14339: out <= 16'hFC97;
    16'd14340: out <= 16'h046E;    16'd14341: out <= 16'h08DC;    16'd14342: out <= 16'hFD0F;    16'd14343: out <= 16'hFEC3;
    16'd14344: out <= 16'hF7E8;    16'd14345: out <= 16'hF9E8;    16'd14346: out <= 16'h0513;    16'd14347: out <= 16'hFD09;
    16'd14348: out <= 16'h01AF;    16'd14349: out <= 16'hFB6A;    16'd14350: out <= 16'hFCAB;    16'd14351: out <= 16'hFD70;
    16'd14352: out <= 16'hFF6C;    16'd14353: out <= 16'h0288;    16'd14354: out <= 16'hFFEF;    16'd14355: out <= 16'h00E9;
    16'd14356: out <= 16'h0383;    16'd14357: out <= 16'h0161;    16'd14358: out <= 16'hFEC8;    16'd14359: out <= 16'hFD4A;
    16'd14360: out <= 16'hFEF6;    16'd14361: out <= 16'hF6E2;    16'd14362: out <= 16'h0388;    16'd14363: out <= 16'h030F;
    16'd14364: out <= 16'hFC8C;    16'd14365: out <= 16'h01B6;    16'd14366: out <= 16'hFF34;    16'd14367: out <= 16'h0239;
    16'd14368: out <= 16'hFE45;    16'd14369: out <= 16'h011D;    16'd14370: out <= 16'h07E2;    16'd14371: out <= 16'h04C6;
    16'd14372: out <= 16'h050A;    16'd14373: out <= 16'h06B2;    16'd14374: out <= 16'h007D;    16'd14375: out <= 16'h03A0;
    16'd14376: out <= 16'h0010;    16'd14377: out <= 16'h008E;    16'd14378: out <= 16'h0023;    16'd14379: out <= 16'h070C;
    16'd14380: out <= 16'hFD1D;    16'd14381: out <= 16'h03D5;    16'd14382: out <= 16'h0A10;    16'd14383: out <= 16'h0818;
    16'd14384: out <= 16'h0102;    16'd14385: out <= 16'h077F;    16'd14386: out <= 16'h0545;    16'd14387: out <= 16'hFBDF;
    16'd14388: out <= 16'hFF85;    16'd14389: out <= 16'h04CE;    16'd14390: out <= 16'h04E6;    16'd14391: out <= 16'h03CC;
    16'd14392: out <= 16'h07D2;    16'd14393: out <= 16'h0156;    16'd14394: out <= 16'h01D8;    16'd14395: out <= 16'h0599;
    16'd14396: out <= 16'h0A0B;    16'd14397: out <= 16'hFF73;    16'd14398: out <= 16'h06E0;    16'd14399: out <= 16'h07AE;
    16'd14400: out <= 16'hFFB0;    16'd14401: out <= 16'h070E;    16'd14402: out <= 16'h034A;    16'd14403: out <= 16'h02BA;
    16'd14404: out <= 16'h04E3;    16'd14405: out <= 16'h00E1;    16'd14406: out <= 16'h05E6;    16'd14407: out <= 16'h07C3;
    16'd14408: out <= 16'h0445;    16'd14409: out <= 16'h06CD;    16'd14410: out <= 16'h07DB;    16'd14411: out <= 16'h005F;
    16'd14412: out <= 16'h0402;    16'd14413: out <= 16'h060E;    16'd14414: out <= 16'h02AB;    16'd14415: out <= 16'h03DF;
    16'd14416: out <= 16'h0691;    16'd14417: out <= 16'h015C;    16'd14418: out <= 16'h08F3;    16'd14419: out <= 16'h02E7;
    16'd14420: out <= 16'hFEB3;    16'd14421: out <= 16'h04CE;    16'd14422: out <= 16'h06DD;    16'd14423: out <= 16'hFBE0;
    16'd14424: out <= 16'hFDF9;    16'd14425: out <= 16'h04FC;    16'd14426: out <= 16'h088D;    16'd14427: out <= 16'h0297;
    16'd14428: out <= 16'h03E6;    16'd14429: out <= 16'h06C8;    16'd14430: out <= 16'h06A4;    16'd14431: out <= 16'h0863;
    16'd14432: out <= 16'h0172;    16'd14433: out <= 16'h029C;    16'd14434: out <= 16'h0060;    16'd14435: out <= 16'h04C8;
    16'd14436: out <= 16'h0002;    16'd14437: out <= 16'h06BC;    16'd14438: out <= 16'h03E3;    16'd14439: out <= 16'h0C6F;
    16'd14440: out <= 16'h0E4C;    16'd14441: out <= 16'h0940;    16'd14442: out <= 16'h0110;    16'd14443: out <= 16'h07C3;
    16'd14444: out <= 16'h00AF;    16'd14445: out <= 16'hFFF3;    16'd14446: out <= 16'h042B;    16'd14447: out <= 16'h029D;
    16'd14448: out <= 16'hFEBE;    16'd14449: out <= 16'h017F;    16'd14450: out <= 16'h04A1;    16'd14451: out <= 16'h0271;
    16'd14452: out <= 16'hFF78;    16'd14453: out <= 16'h0228;    16'd14454: out <= 16'h02F5;    16'd14455: out <= 16'h0A09;
    16'd14456: out <= 16'h0A7B;    16'd14457: out <= 16'h08A7;    16'd14458: out <= 16'h01B5;    16'd14459: out <= 16'h069A;
    16'd14460: out <= 16'h0875;    16'd14461: out <= 16'h0782;    16'd14462: out <= 16'h05E6;    16'd14463: out <= 16'h0A5C;
    16'd14464: out <= 16'h0033;    16'd14465: out <= 16'h04AE;    16'd14466: out <= 16'h0571;    16'd14467: out <= 16'h035E;
    16'd14468: out <= 16'h0418;    16'd14469: out <= 16'h0045;    16'd14470: out <= 16'h0199;    16'd14471: out <= 16'h01E4;
    16'd14472: out <= 16'h064A;    16'd14473: out <= 16'h01E8;    16'd14474: out <= 16'h03E4;    16'd14475: out <= 16'h00B3;
    16'd14476: out <= 16'h01A1;    16'd14477: out <= 16'h0317;    16'd14478: out <= 16'h0143;    16'd14479: out <= 16'h04D9;
    16'd14480: out <= 16'h07FF;    16'd14481: out <= 16'h01A6;    16'd14482: out <= 16'h0424;    16'd14483: out <= 16'h0B76;
    16'd14484: out <= 16'h035A;    16'd14485: out <= 16'h0750;    16'd14486: out <= 16'hFFAC;    16'd14487: out <= 16'h01FF;
    16'd14488: out <= 16'h076B;    16'd14489: out <= 16'h0648;    16'd14490: out <= 16'h0567;    16'd14491: out <= 16'h005C;
    16'd14492: out <= 16'h043D;    16'd14493: out <= 16'h035F;    16'd14494: out <= 16'h02C5;    16'd14495: out <= 16'h0326;
    16'd14496: out <= 16'h078E;    16'd14497: out <= 16'h0729;    16'd14498: out <= 16'h020E;    16'd14499: out <= 16'h0162;
    16'd14500: out <= 16'hFE81;    16'd14501: out <= 16'h08B7;    16'd14502: out <= 16'h0741;    16'd14503: out <= 16'h061F;
    16'd14504: out <= 16'hFAC4;    16'd14505: out <= 16'h00E7;    16'd14506: out <= 16'h0456;    16'd14507: out <= 16'h0839;
    16'd14508: out <= 16'h0AB3;    16'd14509: out <= 16'hFEB4;    16'd14510: out <= 16'h066E;    16'd14511: out <= 16'h0752;
    16'd14512: out <= 16'h0770;    16'd14513: out <= 16'h02CD;    16'd14514: out <= 16'h0866;    16'd14515: out <= 16'h01E8;
    16'd14516: out <= 16'h02E8;    16'd14517: out <= 16'h06BC;    16'd14518: out <= 16'h029C;    16'd14519: out <= 16'h06E2;
    16'd14520: out <= 16'h0876;    16'd14521: out <= 16'h06A9;    16'd14522: out <= 16'hFBB9;    16'd14523: out <= 16'h02E6;
    16'd14524: out <= 16'hFED3;    16'd14525: out <= 16'h0036;    16'd14526: out <= 16'h0329;    16'd14527: out <= 16'h0E20;
    16'd14528: out <= 16'h0378;    16'd14529: out <= 16'h0A48;    16'd14530: out <= 16'h030D;    16'd14531: out <= 16'h0574;
    16'd14532: out <= 16'h0405;    16'd14533: out <= 16'h017C;    16'd14534: out <= 16'h0A38;    16'd14535: out <= 16'hFD21;
    16'd14536: out <= 16'h050F;    16'd14537: out <= 16'h0BD8;    16'd14538: out <= 16'h0345;    16'd14539: out <= 16'h04F8;
    16'd14540: out <= 16'h0477;    16'd14541: out <= 16'h014C;    16'd14542: out <= 16'h0112;    16'd14543: out <= 16'h0231;
    16'd14544: out <= 16'h04ED;    16'd14545: out <= 16'h04A3;    16'd14546: out <= 16'hFD90;    16'd14547: out <= 16'h0059;
    16'd14548: out <= 16'h0638;    16'd14549: out <= 16'h0064;    16'd14550: out <= 16'h013F;    16'd14551: out <= 16'hFB1E;
    16'd14552: out <= 16'hFEB3;    16'd14553: out <= 16'hF8EA;    16'd14554: out <= 16'h0285;    16'd14555: out <= 16'h017A;
    16'd14556: out <= 16'h022C;    16'd14557: out <= 16'hFC65;    16'd14558: out <= 16'hFFF6;    16'd14559: out <= 16'h001E;
    16'd14560: out <= 16'hFD38;    16'd14561: out <= 16'h0429;    16'd14562: out <= 16'h00B5;    16'd14563: out <= 16'hFE6E;
    16'd14564: out <= 16'h003F;    16'd14565: out <= 16'h0088;    16'd14566: out <= 16'hFAEF;    16'd14567: out <= 16'h0042;
    16'd14568: out <= 16'h06DF;    16'd14569: out <= 16'h0100;    16'd14570: out <= 16'hFC60;    16'd14571: out <= 16'h0AD3;
    16'd14572: out <= 16'h02B7;    16'd14573: out <= 16'h05C6;    16'd14574: out <= 16'hFE1D;    16'd14575: out <= 16'h0304;
    16'd14576: out <= 16'hFEBC;    16'd14577: out <= 16'h0158;    16'd14578: out <= 16'h04CE;    16'd14579: out <= 16'hFD24;
    16'd14580: out <= 16'h0148;    16'd14581: out <= 16'h05DC;    16'd14582: out <= 16'h0105;    16'd14583: out <= 16'hF992;
    16'd14584: out <= 16'h016A;    16'd14585: out <= 16'hFDFE;    16'd14586: out <= 16'hFFE1;    16'd14587: out <= 16'hFD2C;
    16'd14588: out <= 16'hFA5D;    16'd14589: out <= 16'h005E;    16'd14590: out <= 16'hFBE5;    16'd14591: out <= 16'h018E;
    16'd14592: out <= 16'h0269;    16'd14593: out <= 16'hFD16;    16'd14594: out <= 16'hF7CD;    16'd14595: out <= 16'h04A9;
    16'd14596: out <= 16'h00CB;    16'd14597: out <= 16'hFA68;    16'd14598: out <= 16'hFC54;    16'd14599: out <= 16'hF958;
    16'd14600: out <= 16'h06D2;    16'd14601: out <= 16'hFB7E;    16'd14602: out <= 16'h0544;    16'd14603: out <= 16'hFE3E;
    16'd14604: out <= 16'h00D4;    16'd14605: out <= 16'h0336;    16'd14606: out <= 16'hF736;    16'd14607: out <= 16'hFEDE;
    16'd14608: out <= 16'hFE1F;    16'd14609: out <= 16'hFAD5;    16'd14610: out <= 16'hFBB5;    16'd14611: out <= 16'h0245;
    16'd14612: out <= 16'hFEF3;    16'd14613: out <= 16'hFF4A;    16'd14614: out <= 16'h002B;    16'd14615: out <= 16'h01D5;
    16'd14616: out <= 16'h0136;    16'd14617: out <= 16'h01A4;    16'd14618: out <= 16'hFC25;    16'd14619: out <= 16'hFBAB;
    16'd14620: out <= 16'h04D4;    16'd14621: out <= 16'hFE3A;    16'd14622: out <= 16'hFF57;    16'd14623: out <= 16'h0773;
    16'd14624: out <= 16'h04C3;    16'd14625: out <= 16'hF896;    16'd14626: out <= 16'h0A31;    16'd14627: out <= 16'h01B5;
    16'd14628: out <= 16'h01CD;    16'd14629: out <= 16'h01FD;    16'd14630: out <= 16'h019A;    16'd14631: out <= 16'h027E;
    16'd14632: out <= 16'h006F;    16'd14633: out <= 16'h039A;    16'd14634: out <= 16'h02BF;    16'd14635: out <= 16'h06F1;
    16'd14636: out <= 16'h0669;    16'd14637: out <= 16'h0812;    16'd14638: out <= 16'h0496;    16'd14639: out <= 16'h053C;
    16'd14640: out <= 16'h02D4;    16'd14641: out <= 16'h080A;    16'd14642: out <= 16'h01D0;    16'd14643: out <= 16'h0078;
    16'd14644: out <= 16'h0015;    16'd14645: out <= 16'h0753;    16'd14646: out <= 16'h0865;    16'd14647: out <= 16'h0165;
    16'd14648: out <= 16'h00D6;    16'd14649: out <= 16'h0303;    16'd14650: out <= 16'h0250;    16'd14651: out <= 16'h08B9;
    16'd14652: out <= 16'h001D;    16'd14653: out <= 16'h0263;    16'd14654: out <= 16'h03DE;    16'd14655: out <= 16'hFFD6;
    16'd14656: out <= 16'h0499;    16'd14657: out <= 16'hFFAA;    16'd14658: out <= 16'hFF9E;    16'd14659: out <= 16'h0A64;
    16'd14660: out <= 16'h04DA;    16'd14661: out <= 16'h0235;    16'd14662: out <= 16'h076A;    16'd14663: out <= 16'h017B;
    16'd14664: out <= 16'h00C3;    16'd14665: out <= 16'h05B1;    16'd14666: out <= 16'h07C1;    16'd14667: out <= 16'hFB9E;
    16'd14668: out <= 16'h056F;    16'd14669: out <= 16'hFFC0;    16'd14670: out <= 16'h0A26;    16'd14671: out <= 16'h04D4;
    16'd14672: out <= 16'h0387;    16'd14673: out <= 16'h02F2;    16'd14674: out <= 16'h030E;    16'd14675: out <= 16'h078D;
    16'd14676: out <= 16'h050D;    16'd14677: out <= 16'h0251;    16'd14678: out <= 16'h0382;    16'd14679: out <= 16'h053A;
    16'd14680: out <= 16'h0A14;    16'd14681: out <= 16'h01CE;    16'd14682: out <= 16'h02D1;    16'd14683: out <= 16'h060E;
    16'd14684: out <= 16'h0008;    16'd14685: out <= 16'h0219;    16'd14686: out <= 16'h04D2;    16'd14687: out <= 16'h0D76;
    16'd14688: out <= 16'h0563;    16'd14689: out <= 16'hFF37;    16'd14690: out <= 16'h09B0;    16'd14691: out <= 16'h0398;
    16'd14692: out <= 16'hFFFD;    16'd14693: out <= 16'h03EC;    16'd14694: out <= 16'h02FB;    16'd14695: out <= 16'h00B3;
    16'd14696: out <= 16'h0831;    16'd14697: out <= 16'h034F;    16'd14698: out <= 16'h040A;    16'd14699: out <= 16'h035D;
    16'd14700: out <= 16'h0248;    16'd14701: out <= 16'h069A;    16'd14702: out <= 16'h0586;    16'd14703: out <= 16'h0776;
    16'd14704: out <= 16'h02BB;    16'd14705: out <= 16'h0374;    16'd14706: out <= 16'h0610;    16'd14707: out <= 16'h0352;
    16'd14708: out <= 16'h02C2;    16'd14709: out <= 16'hFBC7;    16'd14710: out <= 16'h04EC;    16'd14711: out <= 16'h094B;
    16'd14712: out <= 16'h08F9;    16'd14713: out <= 16'h05A8;    16'd14714: out <= 16'h0675;    16'd14715: out <= 16'h03A5;
    16'd14716: out <= 16'h067C;    16'd14717: out <= 16'h03BE;    16'd14718: out <= 16'h00BC;    16'd14719: out <= 16'h0922;
    16'd14720: out <= 16'h02BD;    16'd14721: out <= 16'hFF63;    16'd14722: out <= 16'h01B8;    16'd14723: out <= 16'hFB22;
    16'd14724: out <= 16'h0473;    16'd14725: out <= 16'h04C6;    16'd14726: out <= 16'h00FF;    16'd14727: out <= 16'hFF39;
    16'd14728: out <= 16'h0838;    16'd14729: out <= 16'h055E;    16'd14730: out <= 16'h0344;    16'd14731: out <= 16'hFD1A;
    16'd14732: out <= 16'hFE8A;    16'd14733: out <= 16'h0ABD;    16'd14734: out <= 16'h0659;    16'd14735: out <= 16'h05B1;
    16'd14736: out <= 16'h061B;    16'd14737: out <= 16'h05E4;    16'd14738: out <= 16'h0024;    16'd14739: out <= 16'h0574;
    16'd14740: out <= 16'h0902;    16'd14741: out <= 16'hF8A7;    16'd14742: out <= 16'h0640;    16'd14743: out <= 16'h05E4;
    16'd14744: out <= 16'h0402;    16'd14745: out <= 16'h07F2;    16'd14746: out <= 16'h05E7;    16'd14747: out <= 16'h01E2;
    16'd14748: out <= 16'h03BD;    16'd14749: out <= 16'h011F;    16'd14750: out <= 16'h02AF;    16'd14751: out <= 16'h0476;
    16'd14752: out <= 16'h04D7;    16'd14753: out <= 16'h08DE;    16'd14754: out <= 16'h028D;    16'd14755: out <= 16'hFFFD;
    16'd14756: out <= 16'h04A6;    16'd14757: out <= 16'h01A0;    16'd14758: out <= 16'hFEC0;    16'd14759: out <= 16'h08E3;
    16'd14760: out <= 16'h0281;    16'd14761: out <= 16'h0231;    16'd14762: out <= 16'h0684;    16'd14763: out <= 16'h0522;
    16'd14764: out <= 16'hFEFE;    16'd14765: out <= 16'h022F;    16'd14766: out <= 16'h08DE;    16'd14767: out <= 16'h0574;
    16'd14768: out <= 16'h10BD;    16'd14769: out <= 16'hFFFF;    16'd14770: out <= 16'hFFD2;    16'd14771: out <= 16'hFFF8;
    16'd14772: out <= 16'h06E6;    16'd14773: out <= 16'h0DE8;    16'd14774: out <= 16'h04A9;    16'd14775: out <= 16'h0888;
    16'd14776: out <= 16'h0249;    16'd14777: out <= 16'hFE9B;    16'd14778: out <= 16'h00A1;    16'd14779: out <= 16'h0137;
    16'd14780: out <= 16'h03F8;    16'd14781: out <= 16'h09EB;    16'd14782: out <= 16'h083E;    16'd14783: out <= 16'h0573;
    16'd14784: out <= 16'h06F6;    16'd14785: out <= 16'h086E;    16'd14786: out <= 16'h038D;    16'd14787: out <= 16'h0452;
    16'd14788: out <= 16'h03BA;    16'd14789: out <= 16'h0506;    16'd14790: out <= 16'h009B;    16'd14791: out <= 16'h032A;
    16'd14792: out <= 16'h0820;    16'd14793: out <= 16'hFEC6;    16'd14794: out <= 16'h09E8;    16'd14795: out <= 16'h071E;
    16'd14796: out <= 16'hFD66;    16'd14797: out <= 16'h0560;    16'd14798: out <= 16'h04AE;    16'd14799: out <= 16'hFFD6;
    16'd14800: out <= 16'hFF24;    16'd14801: out <= 16'h0590;    16'd14802: out <= 16'h015F;    16'd14803: out <= 16'h04B5;
    16'd14804: out <= 16'h0632;    16'd14805: out <= 16'h013F;    16'd14806: out <= 16'hFE06;    16'd14807: out <= 16'h05D0;
    16'd14808: out <= 16'hFAD3;    16'd14809: out <= 16'h0334;    16'd14810: out <= 16'h0290;    16'd14811: out <= 16'h0008;
    16'd14812: out <= 16'hFBC9;    16'd14813: out <= 16'hFF59;    16'd14814: out <= 16'hFEC2;    16'd14815: out <= 16'h0298;
    16'd14816: out <= 16'hFEA4;    16'd14817: out <= 16'hFE93;    16'd14818: out <= 16'h00FE;    16'd14819: out <= 16'hFCAD;
    16'd14820: out <= 16'hFF0A;    16'd14821: out <= 16'hFE73;    16'd14822: out <= 16'h0465;    16'd14823: out <= 16'hFCDE;
    16'd14824: out <= 16'h006B;    16'd14825: out <= 16'hFBCE;    16'd14826: out <= 16'h00B9;    16'd14827: out <= 16'h00A8;
    16'd14828: out <= 16'hF94E;    16'd14829: out <= 16'hF955;    16'd14830: out <= 16'hFA12;    16'd14831: out <= 16'hFE6E;
    16'd14832: out <= 16'hFFFF;    16'd14833: out <= 16'hFFF0;    16'd14834: out <= 16'h011A;    16'd14835: out <= 16'hFFC3;
    16'd14836: out <= 16'h0690;    16'd14837: out <= 16'hFE0E;    16'd14838: out <= 16'h0638;    16'd14839: out <= 16'h069C;
    16'd14840: out <= 16'h002E;    16'd14841: out <= 16'h0291;    16'd14842: out <= 16'hFFC4;    16'd14843: out <= 16'hF837;
    16'd14844: out <= 16'h0070;    16'd14845: out <= 16'hFEEF;    16'd14846: out <= 16'hFBC3;    16'd14847: out <= 16'h0083;
    16'd14848: out <= 16'h01D7;    16'd14849: out <= 16'hFF41;    16'd14850: out <= 16'hFA80;    16'd14851: out <= 16'hFC78;
    16'd14852: out <= 16'h01CE;    16'd14853: out <= 16'h040B;    16'd14854: out <= 16'h0162;    16'd14855: out <= 16'hFDD0;
    16'd14856: out <= 16'h01DE;    16'd14857: out <= 16'hFC99;    16'd14858: out <= 16'hFAC5;    16'd14859: out <= 16'h00D5;
    16'd14860: out <= 16'hFBCD;    16'd14861: out <= 16'hFD34;    16'd14862: out <= 16'h0159;    16'd14863: out <= 16'hFE6C;
    16'd14864: out <= 16'hFD04;    16'd14865: out <= 16'hFBDE;    16'd14866: out <= 16'h038D;    16'd14867: out <= 16'h034C;
    16'd14868: out <= 16'h0072;    16'd14869: out <= 16'hFCDE;    16'd14870: out <= 16'h0606;    16'd14871: out <= 16'hFF13;
    16'd14872: out <= 16'hFF39;    16'd14873: out <= 16'h0385;    16'd14874: out <= 16'hFA81;    16'd14875: out <= 16'h0194;
    16'd14876: out <= 16'hFF7C;    16'd14877: out <= 16'hFC1E;    16'd14878: out <= 16'hFD84;    16'd14879: out <= 16'h08D2;
    16'd14880: out <= 16'hFADB;    16'd14881: out <= 16'h02EA;    16'd14882: out <= 16'h0352;    16'd14883: out <= 16'h07F4;
    16'd14884: out <= 16'h0019;    16'd14885: out <= 16'h0142;    16'd14886: out <= 16'h076E;    16'd14887: out <= 16'hFFA9;
    16'd14888: out <= 16'h0307;    16'd14889: out <= 16'hFAAD;    16'd14890: out <= 16'h0760;    16'd14891: out <= 16'hFF7B;
    16'd14892: out <= 16'hFC57;    16'd14893: out <= 16'hFEC4;    16'd14894: out <= 16'h014B;    16'd14895: out <= 16'h0311;
    16'd14896: out <= 16'h03D5;    16'd14897: out <= 16'h01F4;    16'd14898: out <= 16'hFD2E;    16'd14899: out <= 16'h085F;
    16'd14900: out <= 16'h018F;    16'd14901: out <= 16'h06FE;    16'd14902: out <= 16'h013B;    16'd14903: out <= 16'h0A68;
    16'd14904: out <= 16'h0283;    16'd14905: out <= 16'h043B;    16'd14906: out <= 16'h077F;    16'd14907: out <= 16'h0841;
    16'd14908: out <= 16'h02F6;    16'd14909: out <= 16'hFEA9;    16'd14910: out <= 16'h02CB;    16'd14911: out <= 16'h0635;
    16'd14912: out <= 16'h0330;    16'd14913: out <= 16'h02A4;    16'd14914: out <= 16'h0127;    16'd14915: out <= 16'h0337;
    16'd14916: out <= 16'hFFE6;    16'd14917: out <= 16'h027B;    16'd14918: out <= 16'h01CA;    16'd14919: out <= 16'h0745;
    16'd14920: out <= 16'h037F;    16'd14921: out <= 16'h02E2;    16'd14922: out <= 16'h04A8;    16'd14923: out <= 16'h0321;
    16'd14924: out <= 16'h0740;    16'd14925: out <= 16'h0372;    16'd14926: out <= 16'h01EA;    16'd14927: out <= 16'h0180;
    16'd14928: out <= 16'h0253;    16'd14929: out <= 16'h06CC;    16'd14930: out <= 16'h06E6;    16'd14931: out <= 16'h0628;
    16'd14932: out <= 16'h0924;    16'd14933: out <= 16'h0701;    16'd14934: out <= 16'h0203;    16'd14935: out <= 16'h02BC;
    16'd14936: out <= 16'h02F4;    16'd14937: out <= 16'h01D5;    16'd14938: out <= 16'h02E6;    16'd14939: out <= 16'h05D3;
    16'd14940: out <= 16'hFF0F;    16'd14941: out <= 16'h0C1D;    16'd14942: out <= 16'hFAA4;    16'd14943: out <= 16'h088E;
    16'd14944: out <= 16'h0464;    16'd14945: out <= 16'h0033;    16'd14946: out <= 16'h064E;    16'd14947: out <= 16'h01A2;
    16'd14948: out <= 16'h01B3;    16'd14949: out <= 16'h0A80;    16'd14950: out <= 16'h0C40;    16'd14951: out <= 16'h0016;
    16'd14952: out <= 16'h005F;    16'd14953: out <= 16'h03EA;    16'd14954: out <= 16'hFE7E;    16'd14955: out <= 16'h05B1;
    16'd14956: out <= 16'hF9FB;    16'd14957: out <= 16'h0210;    16'd14958: out <= 16'h0079;    16'd14959: out <= 16'h01E2;
    16'd14960: out <= 16'h0969;    16'd14961: out <= 16'h0578;    16'd14962: out <= 16'h075C;    16'd14963: out <= 16'hFFC9;
    16'd14964: out <= 16'h0384;    16'd14965: out <= 16'h0313;    16'd14966: out <= 16'h041F;    16'd14967: out <= 16'h02BA;
    16'd14968: out <= 16'hFEF8;    16'd14969: out <= 16'h044F;    16'd14970: out <= 16'h0135;    16'd14971: out <= 16'h0535;
    16'd14972: out <= 16'h08B2;    16'd14973: out <= 16'h02DF;    16'd14974: out <= 16'h03A8;    16'd14975: out <= 16'h0162;
    16'd14976: out <= 16'h0275;    16'd14977: out <= 16'h0383;    16'd14978: out <= 16'h037E;    16'd14979: out <= 16'h012E;
    16'd14980: out <= 16'h06C2;    16'd14981: out <= 16'hFC2F;    16'd14982: out <= 16'h005F;    16'd14983: out <= 16'h01AD;
    16'd14984: out <= 16'h0795;    16'd14985: out <= 16'h018E;    16'd14986: out <= 16'hFFF6;    16'd14987: out <= 16'h02D7;
    16'd14988: out <= 16'h0A11;    16'd14989: out <= 16'h056E;    16'd14990: out <= 16'h06C0;    16'd14991: out <= 16'h0483;
    16'd14992: out <= 16'h08DA;    16'd14993: out <= 16'h017B;    16'd14994: out <= 16'h065F;    16'd14995: out <= 16'h05DF;
    16'd14996: out <= 16'h0423;    16'd14997: out <= 16'hFFD3;    16'd14998: out <= 16'h0923;    16'd14999: out <= 16'h0280;
    16'd15000: out <= 16'h01FA;    16'd15001: out <= 16'h0635;    16'd15002: out <= 16'h0165;    16'd15003: out <= 16'h05E2;
    16'd15004: out <= 16'h066E;    16'd15005: out <= 16'h04D1;    16'd15006: out <= 16'h06D8;    16'd15007: out <= 16'h00E6;
    16'd15008: out <= 16'h04CC;    16'd15009: out <= 16'h04C9;    16'd15010: out <= 16'h06C4;    16'd15011: out <= 16'h04EC;
    16'd15012: out <= 16'h0542;    16'd15013: out <= 16'h02D7;    16'd15014: out <= 16'h008A;    16'd15015: out <= 16'h0029;
    16'd15016: out <= 16'h0C55;    16'd15017: out <= 16'h0533;    16'd15018: out <= 16'h03A2;    16'd15019: out <= 16'h0A25;
    16'd15020: out <= 16'h0655;    16'd15021: out <= 16'h02D5;    16'd15022: out <= 16'hFD47;    16'd15023: out <= 16'h034E;
    16'd15024: out <= 16'h07AF;    16'd15025: out <= 16'hFFAF;    16'd15026: out <= 16'h03DB;    16'd15027: out <= 16'h0406;
    16'd15028: out <= 16'h05B9;    16'd15029: out <= 16'h00A0;    16'd15030: out <= 16'h040A;    16'd15031: out <= 16'h03C3;
    16'd15032: out <= 16'h077A;    16'd15033: out <= 16'hFFD4;    16'd15034: out <= 16'h048E;    16'd15035: out <= 16'h02DA;
    16'd15036: out <= 16'h06C9;    16'd15037: out <= 16'h0702;    16'd15038: out <= 16'hFE53;    16'd15039: out <= 16'h02FF;
    16'd15040: out <= 16'h07C0;    16'd15041: out <= 16'h06B2;    16'd15042: out <= 16'hFFCB;    16'd15043: out <= 16'hFEDA;
    16'd15044: out <= 16'h02D2;    16'd15045: out <= 16'hFF92;    16'd15046: out <= 16'h00E3;    16'd15047: out <= 16'h02AF;
    16'd15048: out <= 16'h0167;    16'd15049: out <= 16'hFE37;    16'd15050: out <= 16'hFE38;    16'd15051: out <= 16'h055D;
    16'd15052: out <= 16'h04CA;    16'd15053: out <= 16'h0515;    16'd15054: out <= 16'h070D;    16'd15055: out <= 16'h01EE;
    16'd15056: out <= 16'h00C9;    16'd15057: out <= 16'h0A51;    16'd15058: out <= 16'h02F7;    16'd15059: out <= 16'h08E4;
    16'd15060: out <= 16'h00E3;    16'd15061: out <= 16'h049D;    16'd15062: out <= 16'h0504;    16'd15063: out <= 16'h07D5;
    16'd15064: out <= 16'hFADC;    16'd15065: out <= 16'h0284;    16'd15066: out <= 16'h04BB;    16'd15067: out <= 16'h028C;
    16'd15068: out <= 16'h0AC8;    16'd15069: out <= 16'hFB0D;    16'd15070: out <= 16'hFF27;    16'd15071: out <= 16'h02F0;
    16'd15072: out <= 16'hFD93;    16'd15073: out <= 16'hFAD6;    16'd15074: out <= 16'hFF6B;    16'd15075: out <= 16'h0287;
    16'd15076: out <= 16'hFFA1;    16'd15077: out <= 16'hFD62;    16'd15078: out <= 16'h004D;    16'd15079: out <= 16'hFE06;
    16'd15080: out <= 16'h0710;    16'd15081: out <= 16'h0138;    16'd15082: out <= 16'hFF70;    16'd15083: out <= 16'hFE05;
    16'd15084: out <= 16'hFC5B;    16'd15085: out <= 16'h0229;    16'd15086: out <= 16'hFFE4;    16'd15087: out <= 16'hFE59;
    16'd15088: out <= 16'hFD69;    16'd15089: out <= 16'h01A9;    16'd15090: out <= 16'h022B;    16'd15091: out <= 16'hFBEB;
    16'd15092: out <= 16'hF989;    16'd15093: out <= 16'h00F1;    16'd15094: out <= 16'h03B8;    16'd15095: out <= 16'h01CB;
    16'd15096: out <= 16'hF9A6;    16'd15097: out <= 16'h0344;    16'd15098: out <= 16'hFEB2;    16'd15099: out <= 16'h0042;
    16'd15100: out <= 16'hFC0C;    16'd15101: out <= 16'hFA89;    16'd15102: out <= 16'hFF8E;    16'd15103: out <= 16'h00D6;
    16'd15104: out <= 16'h0097;    16'd15105: out <= 16'h02E6;    16'd15106: out <= 16'h0100;    16'd15107: out <= 16'hFDDE;
    16'd15108: out <= 16'hF714;    16'd15109: out <= 16'hFF91;    16'd15110: out <= 16'hFF7E;    16'd15111: out <= 16'hFF9F;
    16'd15112: out <= 16'h03B6;    16'd15113: out <= 16'hFE51;    16'd15114: out <= 16'hFE8C;    16'd15115: out <= 16'h01A8;
    16'd15116: out <= 16'hFCBB;    16'd15117: out <= 16'hF897;    16'd15118: out <= 16'h01E6;    16'd15119: out <= 16'h0336;
    16'd15120: out <= 16'h05CA;    16'd15121: out <= 16'h02E7;    16'd15122: out <= 16'h01DA;    16'd15123: out <= 16'hFE2B;
    16'd15124: out <= 16'hFAB6;    16'd15125: out <= 16'hFF0D;    16'd15126: out <= 16'h097C;    16'd15127: out <= 16'h03AB;
    16'd15128: out <= 16'hFBC5;    16'd15129: out <= 16'hFAFD;    16'd15130: out <= 16'h0196;    16'd15131: out <= 16'hFE73;
    16'd15132: out <= 16'hFE56;    16'd15133: out <= 16'hF82F;    16'd15134: out <= 16'h0397;    16'd15135: out <= 16'h018E;
    16'd15136: out <= 16'h01E0;    16'd15137: out <= 16'hFD2F;    16'd15138: out <= 16'h01CC;    16'd15139: out <= 16'h0A87;
    16'd15140: out <= 16'hFFEB;    16'd15141: out <= 16'h08D6;    16'd15142: out <= 16'h0574;    16'd15143: out <= 16'h02D9;
    16'd15144: out <= 16'h045C;    16'd15145: out <= 16'h004A;    16'd15146: out <= 16'h0438;    16'd15147: out <= 16'h0355;
    16'd15148: out <= 16'h02AA;    16'd15149: out <= 16'h07E3;    16'd15150: out <= 16'hFE00;    16'd15151: out <= 16'h04E1;
    16'd15152: out <= 16'h0540;    16'd15153: out <= 16'h0923;    16'd15154: out <= 16'h061C;    16'd15155: out <= 16'hFF9B;
    16'd15156: out <= 16'h00FE;    16'd15157: out <= 16'h0310;    16'd15158: out <= 16'h0F67;    16'd15159: out <= 16'h046F;
    16'd15160: out <= 16'h0720;    16'd15161: out <= 16'h09CC;    16'd15162: out <= 16'hFA62;    16'd15163: out <= 16'h0363;
    16'd15164: out <= 16'h003D;    16'd15165: out <= 16'h05FD;    16'd15166: out <= 16'h08B6;    16'd15167: out <= 16'h0484;
    16'd15168: out <= 16'h0525;    16'd15169: out <= 16'h06F8;    16'd15170: out <= 16'hFF46;    16'd15171: out <= 16'h0332;
    16'd15172: out <= 16'h0675;    16'd15173: out <= 16'h04C0;    16'd15174: out <= 16'hFE97;    16'd15175: out <= 16'h081F;
    16'd15176: out <= 16'h0876;    16'd15177: out <= 16'h07B3;    16'd15178: out <= 16'h082D;    16'd15179: out <= 16'h0654;
    16'd15180: out <= 16'h0461;    16'd15181: out <= 16'h0345;    16'd15182: out <= 16'hFD8D;    16'd15183: out <= 16'hFA50;
    16'd15184: out <= 16'h02D8;    16'd15185: out <= 16'h0887;    16'd15186: out <= 16'h01BC;    16'd15187: out <= 16'hFF33;
    16'd15188: out <= 16'h0644;    16'd15189: out <= 16'h0442;    16'd15190: out <= 16'h00EA;    16'd15191: out <= 16'h0287;
    16'd15192: out <= 16'h0768;    16'd15193: out <= 16'h03E1;    16'd15194: out <= 16'h0813;    16'd15195: out <= 16'h04DC;
    16'd15196: out <= 16'hFE68;    16'd15197: out <= 16'h02EB;    16'd15198: out <= 16'hFDAD;    16'd15199: out <= 16'h0787;
    16'd15200: out <= 16'h02A5;    16'd15201: out <= 16'h0461;    16'd15202: out <= 16'h048B;    16'd15203: out <= 16'h04C5;
    16'd15204: out <= 16'hFFCC;    16'd15205: out <= 16'h06BA;    16'd15206: out <= 16'hFF59;    16'd15207: out <= 16'h054C;
    16'd15208: out <= 16'h043A;    16'd15209: out <= 16'hFF01;    16'd15210: out <= 16'h0032;    16'd15211: out <= 16'h0454;
    16'd15212: out <= 16'h039E;    16'd15213: out <= 16'h0652;    16'd15214: out <= 16'h0542;    16'd15215: out <= 16'hFE79;
    16'd15216: out <= 16'h0505;    16'd15217: out <= 16'h03AA;    16'd15218: out <= 16'hFE1D;    16'd15219: out <= 16'h0320;
    16'd15220: out <= 16'h05BB;    16'd15221: out <= 16'h06D4;    16'd15222: out <= 16'h01BF;    16'd15223: out <= 16'h041D;
    16'd15224: out <= 16'h096D;    16'd15225: out <= 16'h0016;    16'd15226: out <= 16'hFF15;    16'd15227: out <= 16'h0A2B;
    16'd15228: out <= 16'h0021;    16'd15229: out <= 16'h079A;    16'd15230: out <= 16'h04B5;    16'd15231: out <= 16'h07EE;
    16'd15232: out <= 16'h06E1;    16'd15233: out <= 16'h02B0;    16'd15234: out <= 16'h00D7;    16'd15235: out <= 16'hFDDB;
    16'd15236: out <= 16'h0AA2;    16'd15237: out <= 16'h0549;    16'd15238: out <= 16'h0000;    16'd15239: out <= 16'h0563;
    16'd15240: out <= 16'h05AC;    16'd15241: out <= 16'h06AF;    16'd15242: out <= 16'h0306;    16'd15243: out <= 16'h012C;
    16'd15244: out <= 16'h06C9;    16'd15245: out <= 16'h06BB;    16'd15246: out <= 16'hFCC3;    16'd15247: out <= 16'h06D3;
    16'd15248: out <= 16'h04F1;    16'd15249: out <= 16'hFEA4;    16'd15250: out <= 16'h02C2;    16'd15251: out <= 16'h0169;
    16'd15252: out <= 16'h0208;    16'd15253: out <= 16'h045C;    16'd15254: out <= 16'h0315;    16'd15255: out <= 16'h00B2;
    16'd15256: out <= 16'h0589;    16'd15257: out <= 16'h02BE;    16'd15258: out <= 16'h0061;    16'd15259: out <= 16'h02D3;
    16'd15260: out <= 16'h03BE;    16'd15261: out <= 16'h02C4;    16'd15262: out <= 16'h0298;    16'd15263: out <= 16'h0924;
    16'd15264: out <= 16'h0597;    16'd15265: out <= 16'h0B3C;    16'd15266: out <= 16'h06C5;    16'd15267: out <= 16'h0251;
    16'd15268: out <= 16'h00CA;    16'd15269: out <= 16'h068E;    16'd15270: out <= 16'h09FA;    16'd15271: out <= 16'h012F;
    16'd15272: out <= 16'h076C;    16'd15273: out <= 16'h018C;    16'd15274: out <= 16'h04FF;    16'd15275: out <= 16'hFC79;
    16'd15276: out <= 16'hFDA7;    16'd15277: out <= 16'hFEB2;    16'd15278: out <= 16'h05CF;    16'd15279: out <= 16'h0230;
    16'd15280: out <= 16'hFDF3;    16'd15281: out <= 16'hFEDE;    16'd15282: out <= 16'h04D8;    16'd15283: out <= 16'hFE6A;
    16'd15284: out <= 16'h0332;    16'd15285: out <= 16'h03E0;    16'd15286: out <= 16'h01A4;    16'd15287: out <= 16'h03E0;
    16'd15288: out <= 16'h077B;    16'd15289: out <= 16'h0922;    16'd15290: out <= 16'hFE81;    16'd15291: out <= 16'h0BA8;
    16'd15292: out <= 16'h0BA4;    16'd15293: out <= 16'h051A;    16'd15294: out <= 16'hFF17;    16'd15295: out <= 16'h0136;
    16'd15296: out <= 16'h0015;    16'd15297: out <= 16'h027C;    16'd15298: out <= 16'h0084;    16'd15299: out <= 16'hFC19;
    16'd15300: out <= 16'h05FF;    16'd15301: out <= 16'h0101;    16'd15302: out <= 16'h070B;    16'd15303: out <= 16'hFD5F;
    16'd15304: out <= 16'h0323;    16'd15305: out <= 16'h03C8;    16'd15306: out <= 16'h072D;    16'd15307: out <= 16'hFEDE;
    16'd15308: out <= 16'h05DA;    16'd15309: out <= 16'h047B;    16'd15310: out <= 16'h05CD;    16'd15311: out <= 16'hFFA3;
    16'd15312: out <= 16'h0827;    16'd15313: out <= 16'h08E2;    16'd15314: out <= 16'h03F6;    16'd15315: out <= 16'h02B8;
    16'd15316: out <= 16'h0568;    16'd15317: out <= 16'h0A89;    16'd15318: out <= 16'h08C7;    16'd15319: out <= 16'h01A2;
    16'd15320: out <= 16'hFE5E;    16'd15321: out <= 16'h0589;    16'd15322: out <= 16'hFE94;    16'd15323: out <= 16'hFAF7;
    16'd15324: out <= 16'hFF98;    16'd15325: out <= 16'hFB83;    16'd15326: out <= 16'h01B8;    16'd15327: out <= 16'hFB6C;
    16'd15328: out <= 16'hFBD0;    16'd15329: out <= 16'hFEDC;    16'd15330: out <= 16'hFFCF;    16'd15331: out <= 16'hFA2E;
    16'd15332: out <= 16'hFF35;    16'd15333: out <= 16'h007C;    16'd15334: out <= 16'hFDD5;    16'd15335: out <= 16'h0445;
    16'd15336: out <= 16'hFF24;    16'd15337: out <= 16'hF8D4;    16'd15338: out <= 16'hFB53;    16'd15339: out <= 16'hFE52;
    16'd15340: out <= 16'h0594;    16'd15341: out <= 16'hFDED;    16'd15342: out <= 16'h058C;    16'd15343: out <= 16'hFE92;
    16'd15344: out <= 16'hFDF6;    16'd15345: out <= 16'hFEAA;    16'd15346: out <= 16'hFC09;    16'd15347: out <= 16'h02A8;
    16'd15348: out <= 16'h03E4;    16'd15349: out <= 16'h01AB;    16'd15350: out <= 16'hFC56;    16'd15351: out <= 16'hF950;
    16'd15352: out <= 16'hFF1F;    16'd15353: out <= 16'hFEAC;    16'd15354: out <= 16'hF8BF;    16'd15355: out <= 16'hFDA0;
    16'd15356: out <= 16'hFFA8;    16'd15357: out <= 16'h0333;    16'd15358: out <= 16'h0B3E;    16'd15359: out <= 16'h0009;
    16'd15360: out <= 16'hF923;    16'd15361: out <= 16'h020B;    16'd15362: out <= 16'hFB71;    16'd15363: out <= 16'hFF09;
    16'd15364: out <= 16'hFAAF;    16'd15365: out <= 16'h0067;    16'd15366: out <= 16'h0409;    16'd15367: out <= 16'hF76A;
    16'd15368: out <= 16'h0323;    16'd15369: out <= 16'hFFD6;    16'd15370: out <= 16'h0387;    16'd15371: out <= 16'hFFC4;
    16'd15372: out <= 16'h02A2;    16'd15373: out <= 16'hF95A;    16'd15374: out <= 16'hFF00;    16'd15375: out <= 16'hFF15;
    16'd15376: out <= 16'h0104;    16'd15377: out <= 16'h0046;    16'd15378: out <= 16'h08F0;    16'd15379: out <= 16'h06CD;
    16'd15380: out <= 16'hFB71;    16'd15381: out <= 16'h014F;    16'd15382: out <= 16'h02BE;    16'd15383: out <= 16'h0062;
    16'd15384: out <= 16'h00D4;    16'd15385: out <= 16'h03C7;    16'd15386: out <= 16'hFB8F;    16'd15387: out <= 16'hFA45;
    16'd15388: out <= 16'h02A9;    16'd15389: out <= 16'h02D7;    16'd15390: out <= 16'h0047;    16'd15391: out <= 16'h03CE;
    16'd15392: out <= 16'h0465;    16'd15393: out <= 16'hFEB7;    16'd15394: out <= 16'hFEFC;    16'd15395: out <= 16'h02B9;
    16'd15396: out <= 16'hFC66;    16'd15397: out <= 16'hFF13;    16'd15398: out <= 16'h03FD;    16'd15399: out <= 16'h04EE;
    16'd15400: out <= 16'h0343;    16'd15401: out <= 16'hFF08;    16'd15402: out <= 16'h02C2;    16'd15403: out <= 16'hFFC7;
    16'd15404: out <= 16'h0533;    16'd15405: out <= 16'h043C;    16'd15406: out <= 16'h08F8;    16'd15407: out <= 16'h0072;
    16'd15408: out <= 16'hFFFB;    16'd15409: out <= 16'h0316;    16'd15410: out <= 16'h05E7;    16'd15411: out <= 16'hFC7E;
    16'd15412: out <= 16'hFD5C;    16'd15413: out <= 16'h0B2A;    16'd15414: out <= 16'h0429;    16'd15415: out <= 16'h0112;
    16'd15416: out <= 16'h0421;    16'd15417: out <= 16'h0572;    16'd15418: out <= 16'h06E0;    16'd15419: out <= 16'h0771;
    16'd15420: out <= 16'h0168;    16'd15421: out <= 16'h04F7;    16'd15422: out <= 16'h03D9;    16'd15423: out <= 16'h09EA;
    16'd15424: out <= 16'h0917;    16'd15425: out <= 16'h0434;    16'd15426: out <= 16'h0606;    16'd15427: out <= 16'h0600;
    16'd15428: out <= 16'h0A2D;    16'd15429: out <= 16'h0846;    16'd15430: out <= 16'hFFDC;    16'd15431: out <= 16'h00F5;
    16'd15432: out <= 16'h0479;    16'd15433: out <= 16'h01CD;    16'd15434: out <= 16'h0997;    16'd15435: out <= 16'hFDC3;
    16'd15436: out <= 16'h0574;    16'd15437: out <= 16'h0287;    16'd15438: out <= 16'hFF19;    16'd15439: out <= 16'hFE04;
    16'd15440: out <= 16'h082F;    16'd15441: out <= 16'hFD7F;    16'd15442: out <= 16'h0154;    16'd15443: out <= 16'h072E;
    16'd15444: out <= 16'h08E9;    16'd15445: out <= 16'h06F2;    16'd15446: out <= 16'h0529;    16'd15447: out <= 16'h03F0;
    16'd15448: out <= 16'h0419;    16'd15449: out <= 16'hFE92;    16'd15450: out <= 16'h02AB;    16'd15451: out <= 16'h05FC;
    16'd15452: out <= 16'h09C4;    16'd15453: out <= 16'h0A81;    16'd15454: out <= 16'h03E4;    16'd15455: out <= 16'h034B;
    16'd15456: out <= 16'h0114;    16'd15457: out <= 16'hFF0E;    16'd15458: out <= 16'h0609;    16'd15459: out <= 16'h00FC;
    16'd15460: out <= 16'h03D6;    16'd15461: out <= 16'h056B;    16'd15462: out <= 16'h0B09;    16'd15463: out <= 16'h021A;
    16'd15464: out <= 16'h0172;    16'd15465: out <= 16'h0699;    16'd15466: out <= 16'hFA56;    16'd15467: out <= 16'h091E;
    16'd15468: out <= 16'hFF60;    16'd15469: out <= 16'h0295;    16'd15470: out <= 16'h03C7;    16'd15471: out <= 16'h0921;
    16'd15472: out <= 16'hFE68;    16'd15473: out <= 16'h04A5;    16'd15474: out <= 16'h00FD;    16'd15475: out <= 16'h0364;
    16'd15476: out <= 16'hFF17;    16'd15477: out <= 16'h0A41;    16'd15478: out <= 16'h004C;    16'd15479: out <= 16'h0A89;
    16'd15480: out <= 16'h073C;    16'd15481: out <= 16'h0346;    16'd15482: out <= 16'h0012;    16'd15483: out <= 16'h047D;
    16'd15484: out <= 16'h0249;    16'd15485: out <= 16'h0040;    16'd15486: out <= 16'hFF3A;    16'd15487: out <= 16'h0213;
    16'd15488: out <= 16'h053F;    16'd15489: out <= 16'h0A36;    16'd15490: out <= 16'h0AEE;    16'd15491: out <= 16'h027A;
    16'd15492: out <= 16'h0A03;    16'd15493: out <= 16'hFC3A;    16'd15494: out <= 16'h08BB;    16'd15495: out <= 16'h064A;
    16'd15496: out <= 16'h0206;    16'd15497: out <= 16'h0317;    16'd15498: out <= 16'h03F9;    16'd15499: out <= 16'h0491;
    16'd15500: out <= 16'hFCA3;    16'd15501: out <= 16'h0540;    16'd15502: out <= 16'h0589;    16'd15503: out <= 16'h07EF;
    16'd15504: out <= 16'h0459;    16'd15505: out <= 16'h080E;    16'd15506: out <= 16'h07FD;    16'd15507: out <= 16'h04EB;
    16'd15508: out <= 16'h02E2;    16'd15509: out <= 16'h0547;    16'd15510: out <= 16'h02A8;    16'd15511: out <= 16'h0BF8;
    16'd15512: out <= 16'h0A80;    16'd15513: out <= 16'hFE1E;    16'd15514: out <= 16'h0018;    16'd15515: out <= 16'h085A;
    16'd15516: out <= 16'h074B;    16'd15517: out <= 16'h06D7;    16'd15518: out <= 16'h02E4;    16'd15519: out <= 16'hFCAC;
    16'd15520: out <= 16'h0153;    16'd15521: out <= 16'h0095;    16'd15522: out <= 16'h038A;    16'd15523: out <= 16'h0349;
    16'd15524: out <= 16'h05BF;    16'd15525: out <= 16'h0500;    16'd15526: out <= 16'hFFF3;    16'd15527: out <= 16'h0448;
    16'd15528: out <= 16'hFDF7;    16'd15529: out <= 16'h03E0;    16'd15530: out <= 16'h03BD;    16'd15531: out <= 16'h0153;
    16'd15532: out <= 16'h024C;    16'd15533: out <= 16'h01C2;    16'd15534: out <= 16'h02F9;    16'd15535: out <= 16'h08EA;
    16'd15536: out <= 16'h0691;    16'd15537: out <= 16'h03BA;    16'd15538: out <= 16'h0694;    16'd15539: out <= 16'h0745;
    16'd15540: out <= 16'h069E;    16'd15541: out <= 16'h05BD;    16'd15542: out <= 16'h0289;    16'd15543: out <= 16'h0846;
    16'd15544: out <= 16'h036E;    16'd15545: out <= 16'h0284;    16'd15546: out <= 16'h0532;    16'd15547: out <= 16'h07A7;
    16'd15548: out <= 16'hFE23;    16'd15549: out <= 16'h0140;    16'd15550: out <= 16'h05CC;    16'd15551: out <= 16'h03CD;
    16'd15552: out <= 16'h022D;    16'd15553: out <= 16'h01E6;    16'd15554: out <= 16'h093B;    16'd15555: out <= 16'h046D;
    16'd15556: out <= 16'h01C7;    16'd15557: out <= 16'h045A;    16'd15558: out <= 16'hFCD7;    16'd15559: out <= 16'hFFC3;
    16'd15560: out <= 16'h007A;    16'd15561: out <= 16'h0171;    16'd15562: out <= 16'h0B0F;    16'd15563: out <= 16'h0546;
    16'd15564: out <= 16'hFE93;    16'd15565: out <= 16'hFEB2;    16'd15566: out <= 16'h053B;    16'd15567: out <= 16'h0048;
    16'd15568: out <= 16'h008E;    16'd15569: out <= 16'h0816;    16'd15570: out <= 16'h03C4;    16'd15571: out <= 16'h02D0;
    16'd15572: out <= 16'hFCF9;    16'd15573: out <= 16'h06A5;    16'd15574: out <= 16'h03AB;    16'd15575: out <= 16'h0956;
    16'd15576: out <= 16'h0367;    16'd15577: out <= 16'hFB32;    16'd15578: out <= 16'h0477;    16'd15579: out <= 16'h00F6;
    16'd15580: out <= 16'hFEE3;    16'd15581: out <= 16'hFCE4;    16'd15582: out <= 16'h03E1;    16'd15583: out <= 16'hFC3A;
    16'd15584: out <= 16'hFC3F;    16'd15585: out <= 16'hFD49;    16'd15586: out <= 16'h01FE;    16'd15587: out <= 16'h02FC;
    16'd15588: out <= 16'hFFBD;    16'd15589: out <= 16'h0064;    16'd15590: out <= 16'hFEAB;    16'd15591: out <= 16'h0083;
    16'd15592: out <= 16'h0252;    16'd15593: out <= 16'hFF6F;    16'd15594: out <= 16'h0352;    16'd15595: out <= 16'h0AD4;
    16'd15596: out <= 16'hFFB6;    16'd15597: out <= 16'h076A;    16'd15598: out <= 16'h0001;    16'd15599: out <= 16'hFDB0;
    16'd15600: out <= 16'h0709;    16'd15601: out <= 16'h04E9;    16'd15602: out <= 16'h0085;    16'd15603: out <= 16'h03BB;
    16'd15604: out <= 16'h0229;    16'd15605: out <= 16'h05A8;    16'd15606: out <= 16'h03D0;    16'd15607: out <= 16'h0000;
    16'd15608: out <= 16'hFEC6;    16'd15609: out <= 16'hF88F;    16'd15610: out <= 16'h0410;    16'd15611: out <= 16'h0171;
    16'd15612: out <= 16'hFAE5;    16'd15613: out <= 16'hF9F1;    16'd15614: out <= 16'h065D;    16'd15615: out <= 16'h00FE;
    16'd15616: out <= 16'h01DE;    16'd15617: out <= 16'h02FC;    16'd15618: out <= 16'hF97E;    16'd15619: out <= 16'hFD84;
    16'd15620: out <= 16'h0254;    16'd15621: out <= 16'hFE8A;    16'd15622: out <= 16'h00A9;    16'd15623: out <= 16'h0019;
    16'd15624: out <= 16'h0372;    16'd15625: out <= 16'hFE3D;    16'd15626: out <= 16'hFFD2;    16'd15627: out <= 16'hFE0F;
    16'd15628: out <= 16'h01DB;    16'd15629: out <= 16'h011A;    16'd15630: out <= 16'hFBC9;    16'd15631: out <= 16'hFE7F;
    16'd15632: out <= 16'hF7F6;    16'd15633: out <= 16'hF6D6;    16'd15634: out <= 16'hFC07;    16'd15635: out <= 16'hFC47;
    16'd15636: out <= 16'hFFA7;    16'd15637: out <= 16'h032D;    16'd15638: out <= 16'hFB5F;    16'd15639: out <= 16'hF737;
    16'd15640: out <= 16'hFDD2;    16'd15641: out <= 16'h0134;    16'd15642: out <= 16'h0283;    16'd15643: out <= 16'h0062;
    16'd15644: out <= 16'h00D1;    16'd15645: out <= 16'hFBEF;    16'd15646: out <= 16'hFE4D;    16'd15647: out <= 16'h0544;
    16'd15648: out <= 16'h0F76;    16'd15649: out <= 16'h01C1;    16'd15650: out <= 16'h060E;    16'd15651: out <= 16'h0955;
    16'd15652: out <= 16'h019E;    16'd15653: out <= 16'h026A;    16'd15654: out <= 16'h01CA;    16'd15655: out <= 16'h0450;
    16'd15656: out <= 16'h01C1;    16'd15657: out <= 16'h033A;    16'd15658: out <= 16'h0A3E;    16'd15659: out <= 16'h07BA;
    16'd15660: out <= 16'h05F6;    16'd15661: out <= 16'h0103;    16'd15662: out <= 16'h05CC;    16'd15663: out <= 16'h0322;
    16'd15664: out <= 16'h012F;    16'd15665: out <= 16'h046B;    16'd15666: out <= 16'h0145;    16'd15667: out <= 16'h0424;
    16'd15668: out <= 16'h0451;    16'd15669: out <= 16'h055A;    16'd15670: out <= 16'h0535;    16'd15671: out <= 16'hFB37;
    16'd15672: out <= 16'h08A7;    16'd15673: out <= 16'h0532;    16'd15674: out <= 16'hFCFA;    16'd15675: out <= 16'h04C8;
    16'd15676: out <= 16'h0534;    16'd15677: out <= 16'h069F;    16'd15678: out <= 16'h0606;    16'd15679: out <= 16'h04DD;
    16'd15680: out <= 16'h0025;    16'd15681: out <= 16'h035B;    16'd15682: out <= 16'h04F1;    16'd15683: out <= 16'h0368;
    16'd15684: out <= 16'h0339;    16'd15685: out <= 16'h00C3;    16'd15686: out <= 16'hFFCF;    16'd15687: out <= 16'h0032;
    16'd15688: out <= 16'hFDBE;    16'd15689: out <= 16'h04E8;    16'd15690: out <= 16'h019E;    16'd15691: out <= 16'h03EC;
    16'd15692: out <= 16'h074C;    16'd15693: out <= 16'hFD41;    16'd15694: out <= 16'h0B31;    16'd15695: out <= 16'h04BF;
    16'd15696: out <= 16'h0863;    16'd15697: out <= 16'h011B;    16'd15698: out <= 16'h064D;    16'd15699: out <= 16'h0845;
    16'd15700: out <= 16'h0028;    16'd15701: out <= 16'hFED4;    16'd15702: out <= 16'h061A;    16'd15703: out <= 16'hFC70;
    16'd15704: out <= 16'h0121;    16'd15705: out <= 16'hFEF8;    16'd15706: out <= 16'h0502;    16'd15707: out <= 16'h047A;
    16'd15708: out <= 16'hFD6F;    16'd15709: out <= 16'h001B;    16'd15710: out <= 16'h0605;    16'd15711: out <= 16'h006E;
    16'd15712: out <= 16'h0323;    16'd15713: out <= 16'h00AB;    16'd15714: out <= 16'hFE60;    16'd15715: out <= 16'h0818;
    16'd15716: out <= 16'h0696;    16'd15717: out <= 16'h03AC;    16'd15718: out <= 16'h061E;    16'd15719: out <= 16'h054F;
    16'd15720: out <= 16'h01C4;    16'd15721: out <= 16'hFCCB;    16'd15722: out <= 16'h04CD;    16'd15723: out <= 16'h0A58;
    16'd15724: out <= 16'h0186;    16'd15725: out <= 16'h0414;    16'd15726: out <= 16'h0493;    16'd15727: out <= 16'h021A;
    16'd15728: out <= 16'hFBDC;    16'd15729: out <= 16'h058C;    16'd15730: out <= 16'h03B4;    16'd15731: out <= 16'hFB71;
    16'd15732: out <= 16'h0649;    16'd15733: out <= 16'hFF3C;    16'd15734: out <= 16'h0188;    16'd15735: out <= 16'h00FF;
    16'd15736: out <= 16'h09CE;    16'd15737: out <= 16'h0048;    16'd15738: out <= 16'hFDDE;    16'd15739: out <= 16'h07B6;
    16'd15740: out <= 16'h0606;    16'd15741: out <= 16'h07B4;    16'd15742: out <= 16'h02A0;    16'd15743: out <= 16'h0250;
    16'd15744: out <= 16'h022A;    16'd15745: out <= 16'h0440;    16'd15746: out <= 16'hFE5A;    16'd15747: out <= 16'h02D8;
    16'd15748: out <= 16'hFE9E;    16'd15749: out <= 16'h0448;    16'd15750: out <= 16'h09E8;    16'd15751: out <= 16'h0547;
    16'd15752: out <= 16'h00E2;    16'd15753: out <= 16'h048B;    16'd15754: out <= 16'h01C3;    16'd15755: out <= 16'h0218;
    16'd15756: out <= 16'h040C;    16'd15757: out <= 16'hFE9A;    16'd15758: out <= 16'h0373;    16'd15759: out <= 16'h011D;
    16'd15760: out <= 16'hFDBF;    16'd15761: out <= 16'h0592;    16'd15762: out <= 16'h019C;    16'd15763: out <= 16'h0658;
    16'd15764: out <= 16'h02C3;    16'd15765: out <= 16'h07EF;    16'd15766: out <= 16'h05EA;    16'd15767: out <= 16'h0210;
    16'd15768: out <= 16'h050B;    16'd15769: out <= 16'h046A;    16'd15770: out <= 16'h062C;    16'd15771: out <= 16'h0044;
    16'd15772: out <= 16'h00BF;    16'd15773: out <= 16'hFE37;    16'd15774: out <= 16'h0980;    16'd15775: out <= 16'h0CA9;
    16'd15776: out <= 16'h0326;    16'd15777: out <= 16'h02AA;    16'd15778: out <= 16'h00AD;    16'd15779: out <= 16'h0917;
    16'd15780: out <= 16'h0725;    16'd15781: out <= 16'h045A;    16'd15782: out <= 16'h047F;    16'd15783: out <= 16'h07FD;
    16'd15784: out <= 16'h0373;    16'd15785: out <= 16'h046A;    16'd15786: out <= 16'h06A9;    16'd15787: out <= 16'hFF1E;
    16'd15788: out <= 16'h02B3;    16'd15789: out <= 16'h038F;    16'd15790: out <= 16'h072D;    16'd15791: out <= 16'h0443;
    16'd15792: out <= 16'h00FE;    16'd15793: out <= 16'hFE76;    16'd15794: out <= 16'h01CC;    16'd15795: out <= 16'h03E5;
    16'd15796: out <= 16'h0341;    16'd15797: out <= 16'hFF72;    16'd15798: out <= 16'hFD4F;    16'd15799: out <= 16'h0465;
    16'd15800: out <= 16'h0B19;    16'd15801: out <= 16'h0343;    16'd15802: out <= 16'hFFAB;    16'd15803: out <= 16'h00A5;
    16'd15804: out <= 16'h04B3;    16'd15805: out <= 16'hFFF9;    16'd15806: out <= 16'h04F9;    16'd15807: out <= 16'h0391;
    16'd15808: out <= 16'h066C;    16'd15809: out <= 16'h07A7;    16'd15810: out <= 16'h0947;    16'd15811: out <= 16'h0316;
    16'd15812: out <= 16'h0485;    16'd15813: out <= 16'h05E4;    16'd15814: out <= 16'h0171;    16'd15815: out <= 16'h09F2;
    16'd15816: out <= 16'h0273;    16'd15817: out <= 16'hFE64;    16'd15818: out <= 16'hF942;    16'd15819: out <= 16'h03C7;
    16'd15820: out <= 16'hFCC8;    16'd15821: out <= 16'hFD16;    16'd15822: out <= 16'h03D8;    16'd15823: out <= 16'hFD7A;
    16'd15824: out <= 16'hFB63;    16'd15825: out <= 16'h06FA;    16'd15826: out <= 16'h06B4;    16'd15827: out <= 16'h05B4;
    16'd15828: out <= 16'h04B8;    16'd15829: out <= 16'h022C;    16'd15830: out <= 16'h068A;    16'd15831: out <= 16'h06A4;
    16'd15832: out <= 16'hFC34;    16'd15833: out <= 16'hFFD6;    16'd15834: out <= 16'hFD97;    16'd15835: out <= 16'hFA02;
    16'd15836: out <= 16'h00DA;    16'd15837: out <= 16'hF996;    16'd15838: out <= 16'h0512;    16'd15839: out <= 16'hFE9E;
    16'd15840: out <= 16'hFAE5;    16'd15841: out <= 16'hFF9B;    16'd15842: out <= 16'h00BD;    16'd15843: out <= 16'hFEF2;
    16'd15844: out <= 16'h0196;    16'd15845: out <= 16'hFDEE;    16'd15846: out <= 16'h0600;    16'd15847: out <= 16'hFE4F;
    16'd15848: out <= 16'hFB9D;    16'd15849: out <= 16'h01D7;    16'd15850: out <= 16'h00A8;    16'd15851: out <= 16'hFD05;
    16'd15852: out <= 16'h023D;    16'd15853: out <= 16'hF510;    16'd15854: out <= 16'h02AA;    16'd15855: out <= 16'hFD5E;
    16'd15856: out <= 16'h008F;    16'd15857: out <= 16'h05A3;    16'd15858: out <= 16'hFD0A;    16'd15859: out <= 16'hFA5E;
    16'd15860: out <= 16'h0321;    16'd15861: out <= 16'h0050;    16'd15862: out <= 16'hFEDE;    16'd15863: out <= 16'hFD85;
    16'd15864: out <= 16'h0621;    16'd15865: out <= 16'hFD23;    16'd15866: out <= 16'hFF57;    16'd15867: out <= 16'hFC2A;
    16'd15868: out <= 16'hFB76;    16'd15869: out <= 16'hFA6B;    16'd15870: out <= 16'h075B;    16'd15871: out <= 16'h02D8;
    16'd15872: out <= 16'hFA54;    16'd15873: out <= 16'h0085;    16'd15874: out <= 16'h0374;    16'd15875: out <= 16'hFFE1;
    16'd15876: out <= 16'h0076;    16'd15877: out <= 16'hFD8E;    16'd15878: out <= 16'h0838;    16'd15879: out <= 16'h04F5;
    16'd15880: out <= 16'h0374;    16'd15881: out <= 16'h01E4;    16'd15882: out <= 16'hF47A;    16'd15883: out <= 16'hFBEE;
    16'd15884: out <= 16'h04C7;    16'd15885: out <= 16'h05AA;    16'd15886: out <= 16'hFE8B;    16'd15887: out <= 16'h009F;
    16'd15888: out <= 16'hFD10;    16'd15889: out <= 16'h01B8;    16'd15890: out <= 16'hFC0D;    16'd15891: out <= 16'hFE7F;
    16'd15892: out <= 16'h0113;    16'd15893: out <= 16'hFF85;    16'd15894: out <= 16'hFCD4;    16'd15895: out <= 16'h01E5;
    16'd15896: out <= 16'hFA7E;    16'd15897: out <= 16'h0092;    16'd15898: out <= 16'hFF9D;    16'd15899: out <= 16'hFD51;
    16'd15900: out <= 16'hFBFE;    16'd15901: out <= 16'h051F;    16'd15902: out <= 16'h06CA;    16'd15903: out <= 16'h0A39;
    16'd15904: out <= 16'h0394;    16'd15905: out <= 16'h03BA;    16'd15906: out <= 16'h041B;    16'd15907: out <= 16'h0649;
    16'd15908: out <= 16'h07E4;    16'd15909: out <= 16'h0605;    16'd15910: out <= 16'h0041;    16'd15911: out <= 16'h06F1;
    16'd15912: out <= 16'h01FC;    16'd15913: out <= 16'h0ACF;    16'd15914: out <= 16'h0126;    16'd15915: out <= 16'hFF03;
    16'd15916: out <= 16'h0364;    16'd15917: out <= 16'h05CB;    16'd15918: out <= 16'h070D;    16'd15919: out <= 16'h0389;
    16'd15920: out <= 16'h02B8;    16'd15921: out <= 16'h05A9;    16'd15922: out <= 16'h055C;    16'd15923: out <= 16'h0645;
    16'd15924: out <= 16'h07A8;    16'd15925: out <= 16'h0AC6;    16'd15926: out <= 16'h02D1;    16'd15927: out <= 16'h0ACD;
    16'd15928: out <= 16'h02C9;    16'd15929: out <= 16'hFF0E;    16'd15930: out <= 16'h0790;    16'd15931: out <= 16'h0100;
    16'd15932: out <= 16'h0075;    16'd15933: out <= 16'h0A3A;    16'd15934: out <= 16'h0844;    16'd15935: out <= 16'hFE81;
    16'd15936: out <= 16'h06C2;    16'd15937: out <= 16'h01C6;    16'd15938: out <= 16'h0640;    16'd15939: out <= 16'h0077;
    16'd15940: out <= 16'h0046;    16'd15941: out <= 16'h07F8;    16'd15942: out <= 16'h0537;    16'd15943: out <= 16'h06DC;
    16'd15944: out <= 16'h02D6;    16'd15945: out <= 16'h0A0D;    16'd15946: out <= 16'h00CF;    16'd15947: out <= 16'hFF7A;
    16'd15948: out <= 16'h052D;    16'd15949: out <= 16'h0456;    16'd15950: out <= 16'h0741;    16'd15951: out <= 16'h0612;
    16'd15952: out <= 16'h0AEE;    16'd15953: out <= 16'h050C;    16'd15954: out <= 16'h03B5;    16'd15955: out <= 16'h019C;
    16'd15956: out <= 16'h02EC;    16'd15957: out <= 16'h0485;    16'd15958: out <= 16'h0191;    16'd15959: out <= 16'h04DB;
    16'd15960: out <= 16'hFA76;    16'd15961: out <= 16'hFF32;    16'd15962: out <= 16'h0ABA;    16'd15963: out <= 16'h01C3;
    16'd15964: out <= 16'hFDBD;    16'd15965: out <= 16'h09D2;    16'd15966: out <= 16'hFAFB;    16'd15967: out <= 16'h03B2;
    16'd15968: out <= 16'h05F3;    16'd15969: out <= 16'hF8FB;    16'd15970: out <= 16'hFFF9;    16'd15971: out <= 16'h087E;
    16'd15972: out <= 16'h038F;    16'd15973: out <= 16'h0853;    16'd15974: out <= 16'h0198;    16'd15975: out <= 16'h03B4;
    16'd15976: out <= 16'hFFC3;    16'd15977: out <= 16'h073C;    16'd15978: out <= 16'hFEBC;    16'd15979: out <= 16'h04EC;
    16'd15980: out <= 16'h0A32;    16'd15981: out <= 16'h0443;    16'd15982: out <= 16'hFF68;    16'd15983: out <= 16'h0268;
    16'd15984: out <= 16'h06E0;    16'd15985: out <= 16'h0150;    16'd15986: out <= 16'h0766;    16'd15987: out <= 16'hFF9B;
    16'd15988: out <= 16'h0391;    16'd15989: out <= 16'hFF06;    16'd15990: out <= 16'h0B01;    16'd15991: out <= 16'h005F;
    16'd15992: out <= 16'h07CD;    16'd15993: out <= 16'h0111;    16'd15994: out <= 16'h0505;    16'd15995: out <= 16'h027E;
    16'd15996: out <= 16'h0162;    16'd15997: out <= 16'h02E8;    16'd15998: out <= 16'h073A;    16'd15999: out <= 16'h03DE;
    16'd16000: out <= 16'h078C;    16'd16001: out <= 16'h0617;    16'd16002: out <= 16'h0282;    16'd16003: out <= 16'h0231;
    16'd16004: out <= 16'h0853;    16'd16005: out <= 16'h007F;    16'd16006: out <= 16'hFF67;    16'd16007: out <= 16'h04FC;
    16'd16008: out <= 16'hFA32;    16'd16009: out <= 16'h0964;    16'd16010: out <= 16'h0245;    16'd16011: out <= 16'h06BD;
    16'd16012: out <= 16'h0006;    16'd16013: out <= 16'h002F;    16'd16014: out <= 16'h016B;    16'd16015: out <= 16'h0315;
    16'd16016: out <= 16'h010A;    16'd16017: out <= 16'h054D;    16'd16018: out <= 16'h0A17;    16'd16019: out <= 16'h05CD;
    16'd16020: out <= 16'h02AD;    16'd16021: out <= 16'h07C2;    16'd16022: out <= 16'hFE66;    16'd16023: out <= 16'h0109;
    16'd16024: out <= 16'h0832;    16'd16025: out <= 16'h030C;    16'd16026: out <= 16'h06B9;    16'd16027: out <= 16'h0417;
    16'd16028: out <= 16'hFD42;    16'd16029: out <= 16'h02D5;    16'd16030: out <= 16'h057C;    16'd16031: out <= 16'h02F9;
    16'd16032: out <= 16'hFF85;    16'd16033: out <= 16'h0278;    16'd16034: out <= 16'h0707;    16'd16035: out <= 16'h07FB;
    16'd16036: out <= 16'hFD67;    16'd16037: out <= 16'h0185;    16'd16038: out <= 16'h024D;    16'd16039: out <= 16'h0D8F;
    16'd16040: out <= 16'hFE48;    16'd16041: out <= 16'h0010;    16'd16042: out <= 16'hFE3E;    16'd16043: out <= 16'h03F5;
    16'd16044: out <= 16'h055D;    16'd16045: out <= 16'hFFB6;    16'd16046: out <= 16'h075D;    16'd16047: out <= 16'h0B35;
    16'd16048: out <= 16'h04ED;    16'd16049: out <= 16'h0428;    16'd16050: out <= 16'h040D;    16'd16051: out <= 16'h06B9;
    16'd16052: out <= 16'h05D7;    16'd16053: out <= 16'h00D0;    16'd16054: out <= 16'h00FB;    16'd16055: out <= 16'h0C49;
    16'd16056: out <= 16'hFD36;    16'd16057: out <= 16'h04FE;    16'd16058: out <= 16'h0130;    16'd16059: out <= 16'h051A;
    16'd16060: out <= 16'h02C6;    16'd16061: out <= 16'hFEB4;    16'd16062: out <= 16'h051A;    16'd16063: out <= 16'h0B9C;
    16'd16064: out <= 16'h060A;    16'd16065: out <= 16'hFF4A;    16'd16066: out <= 16'h014D;    16'd16067: out <= 16'h01EA;
    16'd16068: out <= 16'hFFEE;    16'd16069: out <= 16'hFD0E;    16'd16070: out <= 16'h0271;    16'd16071: out <= 16'h02F7;
    16'd16072: out <= 16'hFE8A;    16'd16073: out <= 16'h093B;    16'd16074: out <= 16'h0418;    16'd16075: out <= 16'h00C3;
    16'd16076: out <= 16'hFE8D;    16'd16077: out <= 16'hFDA0;    16'd16078: out <= 16'h05F4;    16'd16079: out <= 16'hFC1D;
    16'd16080: out <= 16'h0654;    16'd16081: out <= 16'h0A4A;    16'd16082: out <= 16'h0175;    16'd16083: out <= 16'hFC3D;
    16'd16084: out <= 16'hF6E3;    16'd16085: out <= 16'h052E;    16'd16086: out <= 16'h0AF2;    16'd16087: out <= 16'h0114;
    16'd16088: out <= 16'h041D;    16'd16089: out <= 16'hFF1E;    16'd16090: out <= 16'hFD59;    16'd16091: out <= 16'h04E0;
    16'd16092: out <= 16'h018A;    16'd16093: out <= 16'h0135;    16'd16094: out <= 16'h00D8;    16'd16095: out <= 16'hFEF3;
    16'd16096: out <= 16'h02C1;    16'd16097: out <= 16'h02C1;    16'd16098: out <= 16'hFC6E;    16'd16099: out <= 16'h0374;
    16'd16100: out <= 16'hFDC0;    16'd16101: out <= 16'h016B;    16'd16102: out <= 16'h022C;    16'd16103: out <= 16'h002D;
    16'd16104: out <= 16'hFE8C;    16'd16105: out <= 16'h041E;    16'd16106: out <= 16'hFF00;    16'd16107: out <= 16'h0178;
    16'd16108: out <= 16'hFEA5;    16'd16109: out <= 16'h0401;    16'd16110: out <= 16'hF980;    16'd16111: out <= 16'hFFA4;
    16'd16112: out <= 16'hFCF9;    16'd16113: out <= 16'hFD32;    16'd16114: out <= 16'hFB06;    16'd16115: out <= 16'h0065;
    16'd16116: out <= 16'h01F2;    16'd16117: out <= 16'h04B9;    16'd16118: out <= 16'hFFC7;    16'd16119: out <= 16'h0522;
    16'd16120: out <= 16'hFF5A;    16'd16121: out <= 16'h0985;    16'd16122: out <= 16'h03C4;    16'd16123: out <= 16'h0784;
    16'd16124: out <= 16'h0753;    16'd16125: out <= 16'hF99D;    16'd16126: out <= 16'hFCB5;    16'd16127: out <= 16'hFC41;
    16'd16128: out <= 16'hFF50;    16'd16129: out <= 16'hFDFD;    16'd16130: out <= 16'hF98B;    16'd16131: out <= 16'hFF15;
    16'd16132: out <= 16'h00AA;    16'd16133: out <= 16'hFED2;    16'd16134: out <= 16'hFB21;    16'd16135: out <= 16'hFE05;
    16'd16136: out <= 16'hFF73;    16'd16137: out <= 16'hFCF9;    16'd16138: out <= 16'hFE1F;    16'd16139: out <= 16'hFDFC;
    16'd16140: out <= 16'h045A;    16'd16141: out <= 16'hFF33;    16'd16142: out <= 16'h0035;    16'd16143: out <= 16'h0152;
    16'd16144: out <= 16'hFF66;    16'd16145: out <= 16'h00AE;    16'd16146: out <= 16'h0529;    16'd16147: out <= 16'h0333;
    16'd16148: out <= 16'hFF66;    16'd16149: out <= 16'h062A;    16'd16150: out <= 16'hFDA8;    16'd16151: out <= 16'hFF3C;
    16'd16152: out <= 16'hFDE8;    16'd16153: out <= 16'hFE35;    16'd16154: out <= 16'hFCAB;    16'd16155: out <= 16'hFEBE;
    16'd16156: out <= 16'hFD84;    16'd16157: out <= 16'hFEB1;    16'd16158: out <= 16'h048D;    16'd16159: out <= 16'h029D;
    16'd16160: out <= 16'h023F;    16'd16161: out <= 16'h06F6;    16'd16162: out <= 16'h061D;    16'd16163: out <= 16'h0506;
    16'd16164: out <= 16'hFE49;    16'd16165: out <= 16'h01C6;    16'd16166: out <= 16'h0333;    16'd16167: out <= 16'hFF9E;
    16'd16168: out <= 16'h0474;    16'd16169: out <= 16'h038C;    16'd16170: out <= 16'h062F;    16'd16171: out <= 16'h0965;
    16'd16172: out <= 16'hFDB1;    16'd16173: out <= 16'h0625;    16'd16174: out <= 16'h023A;    16'd16175: out <= 16'h040B;
    16'd16176: out <= 16'h01C9;    16'd16177: out <= 16'h0094;    16'd16178: out <= 16'h03F4;    16'd16179: out <= 16'h0378;
    16'd16180: out <= 16'h0AA1;    16'd16181: out <= 16'h08FA;    16'd16182: out <= 16'hFBD1;    16'd16183: out <= 16'hFF69;
    16'd16184: out <= 16'h02AE;    16'd16185: out <= 16'h02ED;    16'd16186: out <= 16'h0099;    16'd16187: out <= 16'h07CA;
    16'd16188: out <= 16'h0537;    16'd16189: out <= 16'h04E2;    16'd16190: out <= 16'h0D7C;    16'd16191: out <= 16'h041E;
    16'd16192: out <= 16'h012D;    16'd16193: out <= 16'h023B;    16'd16194: out <= 16'h02F9;    16'd16195: out <= 16'h07D7;
    16'd16196: out <= 16'h06A2;    16'd16197: out <= 16'h0C04;    16'd16198: out <= 16'h0201;    16'd16199: out <= 16'h027B;
    16'd16200: out <= 16'h057B;    16'd16201: out <= 16'h02CB;    16'd16202: out <= 16'h01BC;    16'd16203: out <= 16'h006D;
    16'd16204: out <= 16'h0395;    16'd16205: out <= 16'h0450;    16'd16206: out <= 16'hFF6F;    16'd16207: out <= 16'h04F1;
    16'd16208: out <= 16'h0490;    16'd16209: out <= 16'hFD06;    16'd16210: out <= 16'h06B1;    16'd16211: out <= 16'h01D0;
    16'd16212: out <= 16'h06BB;    16'd16213: out <= 16'h0222;    16'd16214: out <= 16'h0764;    16'd16215: out <= 16'h0417;
    16'd16216: out <= 16'hFB31;    16'd16217: out <= 16'h029C;    16'd16218: out <= 16'hFB36;    16'd16219: out <= 16'h075A;
    16'd16220: out <= 16'hFFEF;    16'd16221: out <= 16'h066D;    16'd16222: out <= 16'h0523;    16'd16223: out <= 16'h01AD;
    16'd16224: out <= 16'h01C8;    16'd16225: out <= 16'h032D;    16'd16226: out <= 16'h02A3;    16'd16227: out <= 16'h00D0;
    16'd16228: out <= 16'hFE56;    16'd16229: out <= 16'h02A9;    16'd16230: out <= 16'h06CA;    16'd16231: out <= 16'h05A4;
    16'd16232: out <= 16'h0415;    16'd16233: out <= 16'h0670;    16'd16234: out <= 16'h05C2;    16'd16235: out <= 16'h0626;
    16'd16236: out <= 16'h0772;    16'd16237: out <= 16'hFEC9;    16'd16238: out <= 16'h06B9;    16'd16239: out <= 16'h021A;
    16'd16240: out <= 16'h029B;    16'd16241: out <= 16'h02E3;    16'd16242: out <= 16'h0610;    16'd16243: out <= 16'h0350;
    16'd16244: out <= 16'hFAB4;    16'd16245: out <= 16'hFF1E;    16'd16246: out <= 16'h09C0;    16'd16247: out <= 16'h06BE;
    16'd16248: out <= 16'h042E;    16'd16249: out <= 16'h055C;    16'd16250: out <= 16'h0543;    16'd16251: out <= 16'h0828;
    16'd16252: out <= 16'h0516;    16'd16253: out <= 16'h044F;    16'd16254: out <= 16'h06E4;    16'd16255: out <= 16'h04C3;
    16'd16256: out <= 16'h03F7;    16'd16257: out <= 16'h0140;    16'd16258: out <= 16'h02ED;    16'd16259: out <= 16'h03DE;
    16'd16260: out <= 16'h016F;    16'd16261: out <= 16'h085C;    16'd16262: out <= 16'h07F8;    16'd16263: out <= 16'h001D;
    16'd16264: out <= 16'h0079;    16'd16265: out <= 16'h01BD;    16'd16266: out <= 16'hFF16;    16'd16267: out <= 16'h0559;
    16'd16268: out <= 16'h03DA;    16'd16269: out <= 16'h04F3;    16'd16270: out <= 16'h00CD;    16'd16271: out <= 16'hFEDB;
    16'd16272: out <= 16'h0395;    16'd16273: out <= 16'h0045;    16'd16274: out <= 16'h012B;    16'd16275: out <= 16'h0724;
    16'd16276: out <= 16'h03E2;    16'd16277: out <= 16'h0855;    16'd16278: out <= 16'h004B;    16'd16279: out <= 16'h01BA;
    16'd16280: out <= 16'hFF83;    16'd16281: out <= 16'h088C;    16'd16282: out <= 16'h0242;    16'd16283: out <= 16'h015A;
    16'd16284: out <= 16'h0472;    16'd16285: out <= 16'h099D;    16'd16286: out <= 16'h03E4;    16'd16287: out <= 16'h0688;
    16'd16288: out <= 16'h0C66;    16'd16289: out <= 16'h03CB;    16'd16290: out <= 16'h0849;    16'd16291: out <= 16'h069F;
    16'd16292: out <= 16'h0AB0;    16'd16293: out <= 16'hFA25;    16'd16294: out <= 16'h0852;    16'd16295: out <= 16'h0AAA;
    16'd16296: out <= 16'h03F6;    16'd16297: out <= 16'hFF8A;    16'd16298: out <= 16'h0E47;    16'd16299: out <= 16'h0479;
    16'd16300: out <= 16'h0300;    16'd16301: out <= 16'hFFEC;    16'd16302: out <= 16'h0025;    16'd16303: out <= 16'h0191;
    16'd16304: out <= 16'h045F;    16'd16305: out <= 16'h0B0B;    16'd16306: out <= 16'h0306;    16'd16307: out <= 16'hFF0B;
    16'd16308: out <= 16'h08BE;    16'd16309: out <= 16'h009E;    16'd16310: out <= 16'hFFC3;    16'd16311: out <= 16'h04B8;
    16'd16312: out <= 16'h073C;    16'd16313: out <= 16'h03BD;    16'd16314: out <= 16'h03F1;    16'd16315: out <= 16'h0547;
    16'd16316: out <= 16'h0498;    16'd16317: out <= 16'h0222;    16'd16318: out <= 16'h0840;    16'd16319: out <= 16'h027A;
    16'd16320: out <= 16'h072E;    16'd16321: out <= 16'h01CF;    16'd16322: out <= 16'h079F;    16'd16323: out <= 16'h014F;
    16'd16324: out <= 16'hFE53;    16'd16325: out <= 16'hFBA8;    16'd16326: out <= 16'h0407;    16'd16327: out <= 16'h0835;
    16'd16328: out <= 16'h03B4;    16'd16329: out <= 16'h01F9;    16'd16330: out <= 16'h032D;    16'd16331: out <= 16'h0838;
    16'd16332: out <= 16'h0535;    16'd16333: out <= 16'h0648;    16'd16334: out <= 16'h072D;    16'd16335: out <= 16'h01B6;
    16'd16336: out <= 16'h0498;    16'd16337: out <= 16'hFCCE;    16'd16338: out <= 16'h03F0;    16'd16339: out <= 16'h0A70;
    16'd16340: out <= 16'h082F;    16'd16341: out <= 16'h01E0;    16'd16342: out <= 16'h0551;    16'd16343: out <= 16'h0C26;
    16'd16344: out <= 16'h0547;    16'd16345: out <= 16'h0134;    16'd16346: out <= 16'hFDA7;    16'd16347: out <= 16'h0065;
    16'd16348: out <= 16'h036E;    16'd16349: out <= 16'h030B;    16'd16350: out <= 16'h04F9;    16'd16351: out <= 16'h03CB;
    16'd16352: out <= 16'h0434;    16'd16353: out <= 16'h021C;    16'd16354: out <= 16'h054F;    16'd16355: out <= 16'hFA75;
    16'd16356: out <= 16'hFF52;    16'd16357: out <= 16'h02EC;    16'd16358: out <= 16'hFF8C;    16'd16359: out <= 16'h058D;
    16'd16360: out <= 16'hFE71;    16'd16361: out <= 16'hFEF8;    16'd16362: out <= 16'h0248;    16'd16363: out <= 16'h0110;
    16'd16364: out <= 16'h0039;    16'd16365: out <= 16'h01C9;    16'd16366: out <= 16'hFFCD;    16'd16367: out <= 16'h0213;
    16'd16368: out <= 16'hFD8D;    16'd16369: out <= 16'hF9A2;    16'd16370: out <= 16'hFE91;    16'd16371: out <= 16'hFEB2;
    16'd16372: out <= 16'hF967;    16'd16373: out <= 16'hFC9F;    16'd16374: out <= 16'hFE06;    16'd16375: out <= 16'h00A8;
    16'd16376: out <= 16'hFEF6;    16'd16377: out <= 16'hFEB3;    16'd16378: out <= 16'hFFDB;    16'd16379: out <= 16'h0637;
    16'd16380: out <= 16'h0375;    16'd16381: out <= 16'h04D1;    16'd16382: out <= 16'h02A1;    16'd16383: out <= 16'hF979;
    16'd16384: out <= 16'h009D;    16'd16385: out <= 16'hFA82;    16'd16386: out <= 16'hFE9D;    16'd16387: out <= 16'h0270;
    16'd16388: out <= 16'hFFDC;    16'd16389: out <= 16'h06DC;    16'd16390: out <= 16'hFD24;    16'd16391: out <= 16'h0053;
    16'd16392: out <= 16'h024C;    16'd16393: out <= 16'h00B8;    16'd16394: out <= 16'h0328;    16'd16395: out <= 16'hFB1B;
    16'd16396: out <= 16'h016A;    16'd16397: out <= 16'h081F;    16'd16398: out <= 16'hF6F0;    16'd16399: out <= 16'hFEF0;
    16'd16400: out <= 16'h0019;    16'd16401: out <= 16'h027B;    16'd16402: out <= 16'h07E1;    16'd16403: out <= 16'hFA24;
    16'd16404: out <= 16'hFFD2;    16'd16405: out <= 16'hFF2B;    16'd16406: out <= 16'hFC5B;    16'd16407: out <= 16'hFEB7;
    16'd16408: out <= 16'h0186;    16'd16409: out <= 16'hFE54;    16'd16410: out <= 16'hFFFC;    16'd16411: out <= 16'h0245;
    16'd16412: out <= 16'hFD80;    16'd16413: out <= 16'hF763;    16'd16414: out <= 16'h032A;    16'd16415: out <= 16'h07F8;
    16'd16416: out <= 16'h057F;    16'd16417: out <= 16'h030E;    16'd16418: out <= 16'h0811;    16'd16419: out <= 16'h0426;
    16'd16420: out <= 16'hFEEF;    16'd16421: out <= 16'h01E4;    16'd16422: out <= 16'h09D7;    16'd16423: out <= 16'h04B9;
    16'd16424: out <= 16'h06AC;    16'd16425: out <= 16'h0C3F;    16'd16426: out <= 16'h0429;    16'd16427: out <= 16'h0856;
    16'd16428: out <= 16'h0722;    16'd16429: out <= 16'h06EC;    16'd16430: out <= 16'h0281;    16'd16431: out <= 16'h0574;
    16'd16432: out <= 16'h0276;    16'd16433: out <= 16'h092B;    16'd16434: out <= 16'hFFA3;    16'd16435: out <= 16'h02A5;
    16'd16436: out <= 16'h074F;    16'd16437: out <= 16'h011D;    16'd16438: out <= 16'h043A;    16'd16439: out <= 16'h05A4;
    16'd16440: out <= 16'h07A3;    16'd16441: out <= 16'h049F;    16'd16442: out <= 16'h0967;    16'd16443: out <= 16'h0244;
    16'd16444: out <= 16'h0236;    16'd16445: out <= 16'hFF75;    16'd16446: out <= 16'h05DE;    16'd16447: out <= 16'h0758;
    16'd16448: out <= 16'h024B;    16'd16449: out <= 16'h088E;    16'd16450: out <= 16'h04AE;    16'd16451: out <= 16'h0188;
    16'd16452: out <= 16'h022E;    16'd16453: out <= 16'h02C3;    16'd16454: out <= 16'h0B54;    16'd16455: out <= 16'h00F6;
    16'd16456: out <= 16'h037D;    16'd16457: out <= 16'h0942;    16'd16458: out <= 16'h01E8;    16'd16459: out <= 16'hFA04;
    16'd16460: out <= 16'h0A4E;    16'd16461: out <= 16'h0027;    16'd16462: out <= 16'h0374;    16'd16463: out <= 16'h090C;
    16'd16464: out <= 16'h004C;    16'd16465: out <= 16'h0882;    16'd16466: out <= 16'h09AF;    16'd16467: out <= 16'h040B;
    16'd16468: out <= 16'h00D4;    16'd16469: out <= 16'hFE28;    16'd16470: out <= 16'hFFD8;    16'd16471: out <= 16'h0389;
    16'd16472: out <= 16'h057B;    16'd16473: out <= 16'h037B;    16'd16474: out <= 16'h07A3;    16'd16475: out <= 16'h04CD;
    16'd16476: out <= 16'h01C5;    16'd16477: out <= 16'h05AB;    16'd16478: out <= 16'h043F;    16'd16479: out <= 16'h09CD;
    16'd16480: out <= 16'h03CC;    16'd16481: out <= 16'h00C1;    16'd16482: out <= 16'h0377;    16'd16483: out <= 16'h01E2;
    16'd16484: out <= 16'h0812;    16'd16485: out <= 16'hFE91;    16'd16486: out <= 16'h0288;    16'd16487: out <= 16'h0079;
    16'd16488: out <= 16'h057E;    16'd16489: out <= 16'h0268;    16'd16490: out <= 16'hFF38;    16'd16491: out <= 16'h0709;
    16'd16492: out <= 16'hFF86;    16'd16493: out <= 16'h07DC;    16'd16494: out <= 16'hFF55;    16'd16495: out <= 16'h09ED;
    16'd16496: out <= 16'h0126;    16'd16497: out <= 16'h04D5;    16'd16498: out <= 16'h02B2;    16'd16499: out <= 16'h0714;
    16'd16500: out <= 16'hFD40;    16'd16501: out <= 16'h07D2;    16'd16502: out <= 16'h0550;    16'd16503: out <= 16'h05B3;
    16'd16504: out <= 16'h0508;    16'd16505: out <= 16'h009D;    16'd16506: out <= 16'h0180;    16'd16507: out <= 16'h04EC;
    16'd16508: out <= 16'h043F;    16'd16509: out <= 16'h0245;    16'd16510: out <= 16'h000C;    16'd16511: out <= 16'h06D5;
    16'd16512: out <= 16'h025E;    16'd16513: out <= 16'h0090;    16'd16514: out <= 16'h04DC;    16'd16515: out <= 16'h01F0;
    16'd16516: out <= 16'h0722;    16'd16517: out <= 16'h0B11;    16'd16518: out <= 16'h08E0;    16'd16519: out <= 16'h048A;
    16'd16520: out <= 16'h07DF;    16'd16521: out <= 16'h0AB5;    16'd16522: out <= 16'hFE6C;    16'd16523: out <= 16'h05B9;
    16'd16524: out <= 16'h0801;    16'd16525: out <= 16'h051E;    16'd16526: out <= 16'h0036;    16'd16527: out <= 16'h0649;
    16'd16528: out <= 16'h0B86;    16'd16529: out <= 16'h03C9;    16'd16530: out <= 16'h0673;    16'd16531: out <= 16'h05F1;
    16'd16532: out <= 16'h0720;    16'd16533: out <= 16'h0871;    16'd16534: out <= 16'h05DA;    16'd16535: out <= 16'h042E;
    16'd16536: out <= 16'h03FB;    16'd16537: out <= 16'h0413;    16'd16538: out <= 16'h0557;    16'd16539: out <= 16'hFDA0;
    16'd16540: out <= 16'h00AE;    16'd16541: out <= 16'h0387;    16'd16542: out <= 16'h069B;    16'd16543: out <= 16'h0528;
    16'd16544: out <= 16'h06BD;    16'd16545: out <= 16'h0427;    16'd16546: out <= 16'h0374;    16'd16547: out <= 16'hFFEF;
    16'd16548: out <= 16'hFF89;    16'd16549: out <= 16'h097B;    16'd16550: out <= 16'h039F;    16'd16551: out <= 16'h03D0;
    16'd16552: out <= 16'h0687;    16'd16553: out <= 16'h02EF;    16'd16554: out <= 16'h02AD;    16'd16555: out <= 16'h001C;
    16'd16556: out <= 16'h013F;    16'd16557: out <= 16'h0555;    16'd16558: out <= 16'hFC84;    16'd16559: out <= 16'h0B0A;
    16'd16560: out <= 16'h08D8;    16'd16561: out <= 16'h0D8B;    16'd16562: out <= 16'h058B;    16'd16563: out <= 16'h017E;
    16'd16564: out <= 16'h05E7;    16'd16565: out <= 16'h018B;    16'd16566: out <= 16'h02ED;    16'd16567: out <= 16'hFF43;
    16'd16568: out <= 16'h02F8;    16'd16569: out <= 16'h07B0;    16'd16570: out <= 16'hFE3D;    16'd16571: out <= 16'hFE93;
    16'd16572: out <= 16'h0851;    16'd16573: out <= 16'h03DD;    16'd16574: out <= 16'h07EB;    16'd16575: out <= 16'h0152;
    16'd16576: out <= 16'hFE95;    16'd16577: out <= 16'h01AF;    16'd16578: out <= 16'h03A8;    16'd16579: out <= 16'h090C;
    16'd16580: out <= 16'h039F;    16'd16581: out <= 16'hFC7E;    16'd16582: out <= 16'hFF58;    16'd16583: out <= 16'h0267;
    16'd16584: out <= 16'h0101;    16'd16585: out <= 16'h003B;    16'd16586: out <= 16'h0072;    16'd16587: out <= 16'hFE6B;
    16'd16588: out <= 16'h0812;    16'd16589: out <= 16'h0961;    16'd16590: out <= 16'h002B;    16'd16591: out <= 16'h0201;
    16'd16592: out <= 16'h09DA;    16'd16593: out <= 16'h0A92;    16'd16594: out <= 16'h0539;    16'd16595: out <= 16'h0A21;
    16'd16596: out <= 16'h04FB;    16'd16597: out <= 16'hFF9C;    16'd16598: out <= 16'hFE0E;    16'd16599: out <= 16'hFF83;
    16'd16600: out <= 16'h0342;    16'd16601: out <= 16'h0600;    16'd16602: out <= 16'hFFFA;    16'd16603: out <= 16'hFE7B;
    16'd16604: out <= 16'h0848;    16'd16605: out <= 16'h009D;    16'd16606: out <= 16'hFFFB;    16'd16607: out <= 16'h011C;
    16'd16608: out <= 16'h03A6;    16'd16609: out <= 16'hFACD;    16'd16610: out <= 16'hFF74;    16'd16611: out <= 16'h010F;
    16'd16612: out <= 16'hFBD1;    16'd16613: out <= 16'hFA71;    16'd16614: out <= 16'hFE64;    16'd16615: out <= 16'hFCC0;
    16'd16616: out <= 16'hFEC2;    16'd16617: out <= 16'h01AE;    16'd16618: out <= 16'h05DC;    16'd16619: out <= 16'hFF87;
    16'd16620: out <= 16'hFB6C;    16'd16621: out <= 16'hFEA8;    16'd16622: out <= 16'hFEC0;    16'd16623: out <= 16'h0065;
    16'd16624: out <= 16'h01E7;    16'd16625: out <= 16'h04B9;    16'd16626: out <= 16'h0196;    16'd16627: out <= 16'hFCB0;
    16'd16628: out <= 16'hFC4C;    16'd16629: out <= 16'h0550;    16'd16630: out <= 16'hFA00;    16'd16631: out <= 16'hFA36;
    16'd16632: out <= 16'h02B3;    16'd16633: out <= 16'h0359;    16'd16634: out <= 16'hFBD8;    16'd16635: out <= 16'hFEA6;
    16'd16636: out <= 16'h031D;    16'd16637: out <= 16'h016F;    16'd16638: out <= 16'hF95C;    16'd16639: out <= 16'hFA3E;
    16'd16640: out <= 16'h0150;    16'd16641: out <= 16'h0852;    16'd16642: out <= 16'hFE3D;    16'd16643: out <= 16'h0528;
    16'd16644: out <= 16'h052F;    16'd16645: out <= 16'h008D;    16'd16646: out <= 16'h03AC;    16'd16647: out <= 16'hFDD4;
    16'd16648: out <= 16'h04FB;    16'd16649: out <= 16'h02FB;    16'd16650: out <= 16'hF903;    16'd16651: out <= 16'h002F;
    16'd16652: out <= 16'h00DA;    16'd16653: out <= 16'h01D3;    16'd16654: out <= 16'h040A;    16'd16655: out <= 16'hFD5C;
    16'd16656: out <= 16'hF9A1;    16'd16657: out <= 16'hF798;    16'd16658: out <= 16'hFEB6;    16'd16659: out <= 16'h03E7;
    16'd16660: out <= 16'h03FA;    16'd16661: out <= 16'hFD2D;    16'd16662: out <= 16'h0045;    16'd16663: out <= 16'hF9A9;
    16'd16664: out <= 16'hFE77;    16'd16665: out <= 16'h0C66;    16'd16666: out <= 16'h031C;    16'd16667: out <= 16'hFD3F;
    16'd16668: out <= 16'hFDBC;    16'd16669: out <= 16'h0045;    16'd16670: out <= 16'hFC4C;    16'd16671: out <= 16'h011B;
    16'd16672: out <= 16'h05BB;    16'd16673: out <= 16'h05E7;    16'd16674: out <= 16'h01B8;    16'd16675: out <= 16'h013A;
    16'd16676: out <= 16'h0974;    16'd16677: out <= 16'h04AB;    16'd16678: out <= 16'h0C41;    16'd16679: out <= 16'h079C;
    16'd16680: out <= 16'hFD7B;    16'd16681: out <= 16'h053D;    16'd16682: out <= 16'h01C6;    16'd16683: out <= 16'h08F6;
    16'd16684: out <= 16'h0663;    16'd16685: out <= 16'h0773;    16'd16686: out <= 16'hFF49;    16'd16687: out <= 16'h069B;
    16'd16688: out <= 16'h07B9;    16'd16689: out <= 16'h014D;    16'd16690: out <= 16'h0A79;    16'd16691: out <= 16'hFC22;
    16'd16692: out <= 16'h053D;    16'd16693: out <= 16'h037F;    16'd16694: out <= 16'h06B7;    16'd16695: out <= 16'h0A62;
    16'd16696: out <= 16'h0189;    16'd16697: out <= 16'h0D2C;    16'd16698: out <= 16'h03EF;    16'd16699: out <= 16'hFAF3;
    16'd16700: out <= 16'hFE89;    16'd16701: out <= 16'h0AB0;    16'd16702: out <= 16'h021B;    16'd16703: out <= 16'h095D;
    16'd16704: out <= 16'h085F;    16'd16705: out <= 16'hFFB2;    16'd16706: out <= 16'h0827;    16'd16707: out <= 16'h058B;
    16'd16708: out <= 16'hFEF5;    16'd16709: out <= 16'h0244;    16'd16710: out <= 16'h01D9;    16'd16711: out <= 16'h0C45;
    16'd16712: out <= 16'h0185;    16'd16713: out <= 16'h0AC6;    16'd16714: out <= 16'h0915;    16'd16715: out <= 16'h0499;
    16'd16716: out <= 16'h0127;    16'd16717: out <= 16'h0798;    16'd16718: out <= 16'h016A;    16'd16719: out <= 16'h032A;
    16'd16720: out <= 16'h05E0;    16'd16721: out <= 16'h03AF;    16'd16722: out <= 16'h02CD;    16'd16723: out <= 16'h05CA;
    16'd16724: out <= 16'h0147;    16'd16725: out <= 16'h02B3;    16'd16726: out <= 16'h0333;    16'd16727: out <= 16'h0843;
    16'd16728: out <= 16'h0381;    16'd16729: out <= 16'h032F;    16'd16730: out <= 16'h0457;    16'd16731: out <= 16'h00E6;
    16'd16732: out <= 16'h05AA;    16'd16733: out <= 16'h067B;    16'd16734: out <= 16'h039C;    16'd16735: out <= 16'h0171;
    16'd16736: out <= 16'h06C4;    16'd16737: out <= 16'h0634;    16'd16738: out <= 16'h0686;    16'd16739: out <= 16'h06BA;
    16'd16740: out <= 16'h031D;    16'd16741: out <= 16'h0634;    16'd16742: out <= 16'h0A1F;    16'd16743: out <= 16'hFB4D;
    16'd16744: out <= 16'h0455;    16'd16745: out <= 16'h0656;    16'd16746: out <= 16'h05A1;    16'd16747: out <= 16'h06FA;
    16'd16748: out <= 16'h0636;    16'd16749: out <= 16'h0956;    16'd16750: out <= 16'h0B3E;    16'd16751: out <= 16'h073E;
    16'd16752: out <= 16'hFF89;    16'd16753: out <= 16'hFA77;    16'd16754: out <= 16'h0221;    16'd16755: out <= 16'h09D9;
    16'd16756: out <= 16'hFD9A;    16'd16757: out <= 16'h0920;    16'd16758: out <= 16'h0520;    16'd16759: out <= 16'h01B4;
    16'd16760: out <= 16'h05DB;    16'd16761: out <= 16'hFC51;    16'd16762: out <= 16'h072E;    16'd16763: out <= 16'h04E7;
    16'd16764: out <= 16'h0347;    16'd16765: out <= 16'h05AC;    16'd16766: out <= 16'hFC7F;    16'd16767: out <= 16'h086B;
    16'd16768: out <= 16'h0583;    16'd16769: out <= 16'h05DB;    16'd16770: out <= 16'h00C8;    16'd16771: out <= 16'h09E2;
    16'd16772: out <= 16'h0114;    16'd16773: out <= 16'hFF62;    16'd16774: out <= 16'h037F;    16'd16775: out <= 16'h00C0;
    16'd16776: out <= 16'h09D8;    16'd16777: out <= 16'hFF5E;    16'd16778: out <= 16'h04B8;    16'd16779: out <= 16'h049D;
    16'd16780: out <= 16'h0724;    16'd16781: out <= 16'h04DA;    16'd16782: out <= 16'h064E;    16'd16783: out <= 16'hFD66;
    16'd16784: out <= 16'h060E;    16'd16785: out <= 16'h02CE;    16'd16786: out <= 16'hFBEF;    16'd16787: out <= 16'hFD96;
    16'd16788: out <= 16'h0784;    16'd16789: out <= 16'hFCF9;    16'd16790: out <= 16'h0578;    16'd16791: out <= 16'h01E3;
    16'd16792: out <= 16'h079E;    16'd16793: out <= 16'h01C5;    16'd16794: out <= 16'hFE3E;    16'd16795: out <= 16'h04A4;
    16'd16796: out <= 16'h021E;    16'd16797: out <= 16'h0560;    16'd16798: out <= 16'h0612;    16'd16799: out <= 16'h0194;
    16'd16800: out <= 16'h073F;    16'd16801: out <= 16'h06E8;    16'd16802: out <= 16'h0227;    16'd16803: out <= 16'hFFDF;
    16'd16804: out <= 16'h0295;    16'd16805: out <= 16'h0532;    16'd16806: out <= 16'h03D8;    16'd16807: out <= 16'h048D;
    16'd16808: out <= 16'h0406;    16'd16809: out <= 16'h0014;    16'd16810: out <= 16'h0987;    16'd16811: out <= 16'h071E;
    16'd16812: out <= 16'h039E;    16'd16813: out <= 16'h00FF;    16'd16814: out <= 16'h00DF;    16'd16815: out <= 16'h019F;
    16'd16816: out <= 16'h0A97;    16'd16817: out <= 16'h00F4;    16'd16818: out <= 16'h0ABC;    16'd16819: out <= 16'h024A;
    16'd16820: out <= 16'h090A;    16'd16821: out <= 16'h0054;    16'd16822: out <= 16'hFE9B;    16'd16823: out <= 16'h0466;
    16'd16824: out <= 16'h06D9;    16'd16825: out <= 16'h01D9;    16'd16826: out <= 16'h085B;    16'd16827: out <= 16'h0A1B;
    16'd16828: out <= 16'hFFDE;    16'd16829: out <= 16'h04DA;    16'd16830: out <= 16'h0085;    16'd16831: out <= 16'h03FB;
    16'd16832: out <= 16'h0B20;    16'd16833: out <= 16'h04BF;    16'd16834: out <= 16'h03CD;    16'd16835: out <= 16'h0B3D;
    16'd16836: out <= 16'h0144;    16'd16837: out <= 16'h076D;    16'd16838: out <= 16'h0579;    16'd16839: out <= 16'h0526;
    16'd16840: out <= 16'h0227;    16'd16841: out <= 16'h0125;    16'd16842: out <= 16'h0565;    16'd16843: out <= 16'h055E;
    16'd16844: out <= 16'h02BC;    16'd16845: out <= 16'h0426;    16'd16846: out <= 16'h0A72;    16'd16847: out <= 16'h050D;
    16'd16848: out <= 16'h02DD;    16'd16849: out <= 16'h0436;    16'd16850: out <= 16'h017C;    16'd16851: out <= 16'h06EE;
    16'd16852: out <= 16'h00B8;    16'd16853: out <= 16'h03F5;    16'd16854: out <= 16'h061B;    16'd16855: out <= 16'h02D5;
    16'd16856: out <= 16'h0211;    16'd16857: out <= 16'h0423;    16'd16858: out <= 16'hFE22;    16'd16859: out <= 16'h02EC;
    16'd16860: out <= 16'hFDAD;    16'd16861: out <= 16'hFDF7;    16'd16862: out <= 16'hFB2A;    16'd16863: out <= 16'h0A4C;
    16'd16864: out <= 16'h01C4;    16'd16865: out <= 16'h04C1;    16'd16866: out <= 16'hF858;    16'd16867: out <= 16'hFFC2;
    16'd16868: out <= 16'h01FB;    16'd16869: out <= 16'hF91B;    16'd16870: out <= 16'hFDEB;    16'd16871: out <= 16'hFA81;
    16'd16872: out <= 16'hFF35;    16'd16873: out <= 16'hFA88;    16'd16874: out <= 16'hFADD;    16'd16875: out <= 16'h078F;
    16'd16876: out <= 16'hFFC9;    16'd16877: out <= 16'h0499;    16'd16878: out <= 16'h02E6;    16'd16879: out <= 16'h022D;
    16'd16880: out <= 16'hFFC1;    16'd16881: out <= 16'hFE1E;    16'd16882: out <= 16'h0227;    16'd16883: out <= 16'h068C;
    16'd16884: out <= 16'h04BD;    16'd16885: out <= 16'hFB5F;    16'd16886: out <= 16'hF776;    16'd16887: out <= 16'hFD9F;
    16'd16888: out <= 16'hFDB8;    16'd16889: out <= 16'hFB2D;    16'd16890: out <= 16'h09E2;    16'd16891: out <= 16'hFE67;
    16'd16892: out <= 16'hFB84;    16'd16893: out <= 16'hFC43;    16'd16894: out <= 16'h0243;    16'd16895: out <= 16'hFD41;
    16'd16896: out <= 16'hFE01;    16'd16897: out <= 16'hFFC7;    16'd16898: out <= 16'h032C;    16'd16899: out <= 16'hFE5E;
    16'd16900: out <= 16'h029D;    16'd16901: out <= 16'h033E;    16'd16902: out <= 16'h0015;    16'd16903: out <= 16'hFF9A;
    16'd16904: out <= 16'hFEFA;    16'd16905: out <= 16'hFA3B;    16'd16906: out <= 16'hFCDE;    16'd16907: out <= 16'hFD65;
    16'd16908: out <= 16'h0232;    16'd16909: out <= 16'h07E3;    16'd16910: out <= 16'h02FA;    16'd16911: out <= 16'hFB87;
    16'd16912: out <= 16'hFC66;    16'd16913: out <= 16'hFCFD;    16'd16914: out <= 16'h061D;    16'd16915: out <= 16'hFA97;
    16'd16916: out <= 16'hF8FC;    16'd16917: out <= 16'h019C;    16'd16918: out <= 16'h039A;    16'd16919: out <= 16'hFFD4;
    16'd16920: out <= 16'h059B;    16'd16921: out <= 16'h02C2;    16'd16922: out <= 16'h0269;    16'd16923: out <= 16'hFBD8;
    16'd16924: out <= 16'h02E8;    16'd16925: out <= 16'h00AB;    16'd16926: out <= 16'h0888;    16'd16927: out <= 16'h0516;
    16'd16928: out <= 16'h054C;    16'd16929: out <= 16'h02A7;    16'd16930: out <= 16'h0006;    16'd16931: out <= 16'h05D9;
    16'd16932: out <= 16'h06C8;    16'd16933: out <= 16'hFF14;    16'd16934: out <= 16'h0C90;    16'd16935: out <= 16'h0770;
    16'd16936: out <= 16'h0A69;    16'd16937: out <= 16'h04E3;    16'd16938: out <= 16'h044D;    16'd16939: out <= 16'h028E;
    16'd16940: out <= 16'h0006;    16'd16941: out <= 16'h0110;    16'd16942: out <= 16'h058C;    16'd16943: out <= 16'h0123;
    16'd16944: out <= 16'h0420;    16'd16945: out <= 16'hFFDA;    16'd16946: out <= 16'hFCB6;    16'd16947: out <= 16'hFDC3;
    16'd16948: out <= 16'h059E;    16'd16949: out <= 16'h0A24;    16'd16950: out <= 16'h0742;    16'd16951: out <= 16'h0118;
    16'd16952: out <= 16'h05EA;    16'd16953: out <= 16'h0150;    16'd16954: out <= 16'h0579;    16'd16955: out <= 16'hFDC6;
    16'd16956: out <= 16'h05E6;    16'd16957: out <= 16'h073E;    16'd16958: out <= 16'h0881;    16'd16959: out <= 16'h092B;
    16'd16960: out <= 16'h0232;    16'd16961: out <= 16'h0173;    16'd16962: out <= 16'h0655;    16'd16963: out <= 16'h02F3;
    16'd16964: out <= 16'h043F;    16'd16965: out <= 16'h0129;    16'd16966: out <= 16'h00C9;    16'd16967: out <= 16'h04F6;
    16'd16968: out <= 16'hFD6D;    16'd16969: out <= 16'h0648;    16'd16970: out <= 16'h0258;    16'd16971: out <= 16'h0790;
    16'd16972: out <= 16'hFFC9;    16'd16973: out <= 16'h030E;    16'd16974: out <= 16'h04F9;    16'd16975: out <= 16'h0324;
    16'd16976: out <= 16'h041A;    16'd16977: out <= 16'h0A9B;    16'd16978: out <= 16'h0974;    16'd16979: out <= 16'hFF55;
    16'd16980: out <= 16'h069D;    16'd16981: out <= 16'hFF9F;    16'd16982: out <= 16'h05D1;    16'd16983: out <= 16'h06EF;
    16'd16984: out <= 16'h07CD;    16'd16985: out <= 16'h0437;    16'd16986: out <= 16'h0530;    16'd16987: out <= 16'h057F;
    16'd16988: out <= 16'h0328;    16'd16989: out <= 16'hFF4D;    16'd16990: out <= 16'h0395;    16'd16991: out <= 16'h0072;
    16'd16992: out <= 16'hFE45;    16'd16993: out <= 16'h06A7;    16'd16994: out <= 16'h0318;    16'd16995: out <= 16'h044C;
    16'd16996: out <= 16'h02AA;    16'd16997: out <= 16'h0901;    16'd16998: out <= 16'h0315;    16'd16999: out <= 16'h014D;
    16'd17000: out <= 16'h07BB;    16'd17001: out <= 16'h0112;    16'd17002: out <= 16'h06DA;    16'd17003: out <= 16'hFF26;
    16'd17004: out <= 16'h05F0;    16'd17005: out <= 16'h04E6;    16'd17006: out <= 16'h0973;    16'd17007: out <= 16'h064D;
    16'd17008: out <= 16'hFE28;    16'd17009: out <= 16'h03F5;    16'd17010: out <= 16'h072D;    16'd17011: out <= 16'h0168;
    16'd17012: out <= 16'h08D6;    16'd17013: out <= 16'h015F;    16'd17014: out <= 16'hFDC6;    16'd17015: out <= 16'h04F8;
    16'd17016: out <= 16'h0372;    16'd17017: out <= 16'hFDA1;    16'd17018: out <= 16'h0A60;    16'd17019: out <= 16'hFF8F;
    16'd17020: out <= 16'h0390;    16'd17021: out <= 16'h06E7;    16'd17022: out <= 16'h0476;    16'd17023: out <= 16'h08C3;
    16'd17024: out <= 16'h0CDC;    16'd17025: out <= 16'h0706;    16'd17026: out <= 16'h0195;    16'd17027: out <= 16'h0219;
    16'd17028: out <= 16'h02BD;    16'd17029: out <= 16'h02FE;    16'd17030: out <= 16'h0782;    16'd17031: out <= 16'h05E6;
    16'd17032: out <= 16'h0262;    16'd17033: out <= 16'h076A;    16'd17034: out <= 16'hFE95;    16'd17035: out <= 16'h05E7;
    16'd17036: out <= 16'h0888;    16'd17037: out <= 16'h09AB;    16'd17038: out <= 16'h0151;    16'd17039: out <= 16'h04CA;
    16'd17040: out <= 16'h0779;    16'd17041: out <= 16'hFC45;    16'd17042: out <= 16'h09EC;    16'd17043: out <= 16'h071A;
    16'd17044: out <= 16'h096C;    16'd17045: out <= 16'h04A5;    16'd17046: out <= 16'h0267;    16'd17047: out <= 16'h0C4F;
    16'd17048: out <= 16'hFEAE;    16'd17049: out <= 16'h01AB;    16'd17050: out <= 16'h09D5;    16'd17051: out <= 16'h0D1D;
    16'd17052: out <= 16'h0B42;    16'd17053: out <= 16'h061A;    16'd17054: out <= 16'h08C4;    16'd17055: out <= 16'h0357;
    16'd17056: out <= 16'h03B9;    16'd17057: out <= 16'h06E4;    16'd17058: out <= 16'h04C9;    16'd17059: out <= 16'h02A2;
    16'd17060: out <= 16'h0A93;    16'd17061: out <= 16'h0608;    16'd17062: out <= 16'hFD3D;    16'd17063: out <= 16'h016F;
    16'd17064: out <= 16'h0576;    16'd17065: out <= 16'hFF77;    16'd17066: out <= 16'h00BD;    16'd17067: out <= 16'h0AA8;
    16'd17068: out <= 16'hFE44;    16'd17069: out <= 16'h0733;    16'd17070: out <= 16'h0263;    16'd17071: out <= 16'h006B;
    16'd17072: out <= 16'h040F;    16'd17073: out <= 16'h047E;    16'd17074: out <= 16'h0030;    16'd17075: out <= 16'h0204;
    16'd17076: out <= 16'h0AF3;    16'd17077: out <= 16'h097E;    16'd17078: out <= 16'h061F;    16'd17079: out <= 16'h02C2;
    16'd17080: out <= 16'h0C29;    16'd17081: out <= 16'h060E;    16'd17082: out <= 16'hFB3C;    16'd17083: out <= 16'h018D;
    16'd17084: out <= 16'h00D2;    16'd17085: out <= 16'h08EE;    16'd17086: out <= 16'h0552;    16'd17087: out <= 16'h0A1C;
    16'd17088: out <= 16'hFB35;    16'd17089: out <= 16'h07B2;    16'd17090: out <= 16'h0474;    16'd17091: out <= 16'h065B;
    16'd17092: out <= 16'h04E2;    16'd17093: out <= 16'h05F6;    16'd17094: out <= 16'h010C;    16'd17095: out <= 16'h0419;
    16'd17096: out <= 16'h003B;    16'd17097: out <= 16'h02A8;    16'd17098: out <= 16'h025C;    16'd17099: out <= 16'h0866;
    16'd17100: out <= 16'h0A37;    16'd17101: out <= 16'h0258;    16'd17102: out <= 16'h0358;    16'd17103: out <= 16'h04E1;
    16'd17104: out <= 16'h07C8;    16'd17105: out <= 16'h0250;    16'd17106: out <= 16'h04D9;    16'd17107: out <= 16'h07CF;
    16'd17108: out <= 16'h0C81;    16'd17109: out <= 16'h019A;    16'd17110: out <= 16'hFE11;    16'd17111: out <= 16'h04FB;
    16'd17112: out <= 16'h0324;    16'd17113: out <= 16'h06C4;    16'd17114: out <= 16'h025D;    16'd17115: out <= 16'h03A0;
    16'd17116: out <= 16'h00E8;    16'd17117: out <= 16'hFE3F;    16'd17118: out <= 16'hFEC2;    16'd17119: out <= 16'hFF8C;
    16'd17120: out <= 16'hFCC2;    16'd17121: out <= 16'h022D;    16'd17122: out <= 16'h02F8;    16'd17123: out <= 16'h005F;
    16'd17124: out <= 16'hFD08;    16'd17125: out <= 16'hFD71;    16'd17126: out <= 16'h01D4;    16'd17127: out <= 16'hFF82;
    16'd17128: out <= 16'hFBCA;    16'd17129: out <= 16'hFD3E;    16'd17130: out <= 16'h0778;    16'd17131: out <= 16'hFF97;
    16'd17132: out <= 16'hFCCF;    16'd17133: out <= 16'hF9A0;    16'd17134: out <= 16'hFE22;    16'd17135: out <= 16'hFED6;
    16'd17136: out <= 16'h002E;    16'd17137: out <= 16'hFFC3;    16'd17138: out <= 16'hFBAF;    16'd17139: out <= 16'hFCA1;
    16'd17140: out <= 16'hFD3E;    16'd17141: out <= 16'hFBAC;    16'd17142: out <= 16'hFF11;    16'd17143: out <= 16'h03B2;
    16'd17144: out <= 16'h01FB;    16'd17145: out <= 16'hFAF0;    16'd17146: out <= 16'h0ED3;    16'd17147: out <= 16'h02B8;
    16'd17148: out <= 16'h0031;    16'd17149: out <= 16'hF991;    16'd17150: out <= 16'hFFC9;    16'd17151: out <= 16'hFE34;
    16'd17152: out <= 16'hFCE1;    16'd17153: out <= 16'hFAE5;    16'd17154: out <= 16'hFF10;    16'd17155: out <= 16'h01BC;
    16'd17156: out <= 16'h07D7;    16'd17157: out <= 16'h00B9;    16'd17158: out <= 16'h0140;    16'd17159: out <= 16'h01C0;
    16'd17160: out <= 16'h0163;    16'd17161: out <= 16'hFCC4;    16'd17162: out <= 16'h04C1;    16'd17163: out <= 16'hFC2F;
    16'd17164: out <= 16'hFCC3;    16'd17165: out <= 16'hFF1E;    16'd17166: out <= 16'h0268;    16'd17167: out <= 16'hFC32;
    16'd17168: out <= 16'hFD53;    16'd17169: out <= 16'h010A;    16'd17170: out <= 16'h0049;    16'd17171: out <= 16'h01D4;
    16'd17172: out <= 16'hFA07;    16'd17173: out <= 16'h077C;    16'd17174: out <= 16'h0690;    16'd17175: out <= 16'h08F7;
    16'd17176: out <= 16'h07F9;    16'd17177: out <= 16'h00A9;    16'd17178: out <= 16'hFFF4;    16'd17179: out <= 16'h00B1;
    16'd17180: out <= 16'hFE94;    16'd17181: out <= 16'h01BC;    16'd17182: out <= 16'hFB93;    16'd17183: out <= 16'h09A2;
    16'd17184: out <= 16'hFD17;    16'd17185: out <= 16'h00C0;    16'd17186: out <= 16'h07A3;    16'd17187: out <= 16'h03AA;
    16'd17188: out <= 16'h07CC;    16'd17189: out <= 16'hFE92;    16'd17190: out <= 16'h06F6;    16'd17191: out <= 16'h07FA;
    16'd17192: out <= 16'h0493;    16'd17193: out <= 16'hFFE5;    16'd17194: out <= 16'hFF3B;    16'd17195: out <= 16'h0206;
    16'd17196: out <= 16'h072A;    16'd17197: out <= 16'h05F1;    16'd17198: out <= 16'hFDB4;    16'd17199: out <= 16'h0565;
    16'd17200: out <= 16'hFE2A;    16'd17201: out <= 16'h02FF;    16'd17202: out <= 16'h02BF;    16'd17203: out <= 16'h0A57;
    16'd17204: out <= 16'h0214;    16'd17205: out <= 16'hFFC5;    16'd17206: out <= 16'h00D5;    16'd17207: out <= 16'hFDC9;
    16'd17208: out <= 16'hFF09;    16'd17209: out <= 16'h068F;    16'd17210: out <= 16'hFFBD;    16'd17211: out <= 16'h0207;
    16'd17212: out <= 16'h008D;    16'd17213: out <= 16'h04AA;    16'd17214: out <= 16'h066D;    16'd17215: out <= 16'hFF6A;
    16'd17216: out <= 16'h03EC;    16'd17217: out <= 16'h024F;    16'd17218: out <= 16'h08B1;    16'd17219: out <= 16'h0A99;
    16'd17220: out <= 16'h04CD;    16'd17221: out <= 16'h04A6;    16'd17222: out <= 16'h06AE;    16'd17223: out <= 16'h0547;
    16'd17224: out <= 16'hFECA;    16'd17225: out <= 16'h067C;    16'd17226: out <= 16'hFE2D;    16'd17227: out <= 16'h09B5;
    16'd17228: out <= 16'hFF63;    16'd17229: out <= 16'h0016;    16'd17230: out <= 16'h0122;    16'd17231: out <= 16'h0458;
    16'd17232: out <= 16'h0892;    16'd17233: out <= 16'h00AF;    16'd17234: out <= 16'h014E;    16'd17235: out <= 16'h08DB;
    16'd17236: out <= 16'h0493;    16'd17237: out <= 16'h01AE;    16'd17238: out <= 16'h022C;    16'd17239: out <= 16'h074B;
    16'd17240: out <= 16'hFE3C;    16'd17241: out <= 16'h08CE;    16'd17242: out <= 16'h03EF;    16'd17243: out <= 16'hFF84;
    16'd17244: out <= 16'h0840;    16'd17245: out <= 16'h0507;    16'd17246: out <= 16'h0307;    16'd17247: out <= 16'h0142;
    16'd17248: out <= 16'h04D8;    16'd17249: out <= 16'h0247;    16'd17250: out <= 16'h016D;    16'd17251: out <= 16'h064F;
    16'd17252: out <= 16'h072C;    16'd17253: out <= 16'hFE21;    16'd17254: out <= 16'h0C6A;    16'd17255: out <= 16'h0057;
    16'd17256: out <= 16'h06A3;    16'd17257: out <= 16'h0C4F;    16'd17258: out <= 16'h06E8;    16'd17259: out <= 16'h0810;
    16'd17260: out <= 16'h0458;    16'd17261: out <= 16'h08ED;    16'd17262: out <= 16'h097D;    16'd17263: out <= 16'h01A5;
    16'd17264: out <= 16'h05B7;    16'd17265: out <= 16'h0118;    16'd17266: out <= 16'h047E;    16'd17267: out <= 16'h063A;
    16'd17268: out <= 16'h064A;    16'd17269: out <= 16'h05A1;    16'd17270: out <= 16'h05F6;    16'd17271: out <= 16'h06A9;
    16'd17272: out <= 16'h02BC;    16'd17273: out <= 16'h0729;    16'd17274: out <= 16'h0388;    16'd17275: out <= 16'h024B;
    16'd17276: out <= 16'h0A12;    16'd17277: out <= 16'h0245;    16'd17278: out <= 16'h0207;    16'd17279: out <= 16'h05DD;
    16'd17280: out <= 16'hFDB3;    16'd17281: out <= 16'h00E6;    16'd17282: out <= 16'hFAB1;    16'd17283: out <= 16'h066F;
    16'd17284: out <= 16'h03A4;    16'd17285: out <= 16'h06E6;    16'd17286: out <= 16'hFFD0;    16'd17287: out <= 16'h0633;
    16'd17288: out <= 16'hFDE5;    16'd17289: out <= 16'h07BF;    16'd17290: out <= 16'h084F;    16'd17291: out <= 16'h09FE;
    16'd17292: out <= 16'h01C2;    16'd17293: out <= 16'h0969;    16'd17294: out <= 16'h06C6;    16'd17295: out <= 16'h04A1;
    16'd17296: out <= 16'hFE84;    16'd17297: out <= 16'h0A14;    16'd17298: out <= 16'h0A26;    16'd17299: out <= 16'h01F9;
    16'd17300: out <= 16'h08E9;    16'd17301: out <= 16'h0690;    16'd17302: out <= 16'h0739;    16'd17303: out <= 16'h05B6;
    16'd17304: out <= 16'hFF6A;    16'd17305: out <= 16'h058B;    16'd17306: out <= 16'h071B;    16'd17307: out <= 16'h022A;
    16'd17308: out <= 16'h051A;    16'd17309: out <= 16'h00C6;    16'd17310: out <= 16'h01A9;    16'd17311: out <= 16'hFF8B;
    16'd17312: out <= 16'h0401;    16'd17313: out <= 16'h0444;    16'd17314: out <= 16'h097B;    16'd17315: out <= 16'hFD5C;
    16'd17316: out <= 16'h01CE;    16'd17317: out <= 16'h0154;    16'd17318: out <= 16'h0219;    16'd17319: out <= 16'h05AF;
    16'd17320: out <= 16'h0473;    16'd17321: out <= 16'h0277;    16'd17322: out <= 16'h02A6;    16'd17323: out <= 16'h0187;
    16'd17324: out <= 16'h069D;    16'd17325: out <= 16'h0662;    16'd17326: out <= 16'h0549;    16'd17327: out <= 16'h0769;
    16'd17328: out <= 16'hFD16;    16'd17329: out <= 16'h00C7;    16'd17330: out <= 16'h07E3;    16'd17331: out <= 16'h00E6;
    16'd17332: out <= 16'h06C4;    16'd17333: out <= 16'h03D3;    16'd17334: out <= 16'h016F;    16'd17335: out <= 16'h06E4;
    16'd17336: out <= 16'h01C4;    16'd17337: out <= 16'h002B;    16'd17338: out <= 16'h053B;    16'd17339: out <= 16'h0B21;
    16'd17340: out <= 16'h0869;    16'd17341: out <= 16'hFEF5;    16'd17342: out <= 16'h0445;    16'd17343: out <= 16'hFC99;
    16'd17344: out <= 16'h010E;    16'd17345: out <= 16'h0129;    16'd17346: out <= 16'h0350;    16'd17347: out <= 16'h00B8;
    16'd17348: out <= 16'hFE3B;    16'd17349: out <= 16'h098C;    16'd17350: out <= 16'h0141;    16'd17351: out <= 16'h05CB;
    16'd17352: out <= 16'h07D6;    16'd17353: out <= 16'h01D2;    16'd17354: out <= 16'h0220;    16'd17355: out <= 16'h09A5;
    16'd17356: out <= 16'h04F0;    16'd17357: out <= 16'h0E70;    16'd17358: out <= 16'h0377;    16'd17359: out <= 16'h05E6;
    16'd17360: out <= 16'h0502;    16'd17361: out <= 16'h03CF;    16'd17362: out <= 16'h06C4;    16'd17363: out <= 16'h02FE;
    16'd17364: out <= 16'hFE71;    16'd17365: out <= 16'h08C6;    16'd17366: out <= 16'h0874;    16'd17367: out <= 16'h0357;
    16'd17368: out <= 16'h025B;    16'd17369: out <= 16'h02F7;    16'd17370: out <= 16'hFA2B;    16'd17371: out <= 16'hFE84;
    16'd17372: out <= 16'hFF0C;    16'd17373: out <= 16'hFFB7;    16'd17374: out <= 16'h0635;    16'd17375: out <= 16'hFF56;
    16'd17376: out <= 16'hFFE2;    16'd17377: out <= 16'h000D;    16'd17378: out <= 16'hFAF1;    16'd17379: out <= 16'h0242;
    16'd17380: out <= 16'hFFD9;    16'd17381: out <= 16'h078B;    16'd17382: out <= 16'hFB42;    16'd17383: out <= 16'h0005;
    16'd17384: out <= 16'h0135;    16'd17385: out <= 16'hFE67;    16'd17386: out <= 16'hFA43;    16'd17387: out <= 16'h07CB;
    16'd17388: out <= 16'h05D2;    16'd17389: out <= 16'h0086;    16'd17390: out <= 16'hF901;    16'd17391: out <= 16'hFDA0;
    16'd17392: out <= 16'hF9F1;    16'd17393: out <= 16'h007F;    16'd17394: out <= 16'h000E;    16'd17395: out <= 16'h024C;
    16'd17396: out <= 16'hFCEF;    16'd17397: out <= 16'hFF04;    16'd17398: out <= 16'hFE70;    16'd17399: out <= 16'h0447;
    16'd17400: out <= 16'hFF78;    16'd17401: out <= 16'hFE34;    16'd17402: out <= 16'hFE01;    16'd17403: out <= 16'h012C;
    16'd17404: out <= 16'hFC64;    16'd17405: out <= 16'h013C;    16'd17406: out <= 16'h0181;    16'd17407: out <= 16'hFAB8;
    16'd17408: out <= 16'h061A;    16'd17409: out <= 16'h057E;    16'd17410: out <= 16'hFDA6;    16'd17411: out <= 16'hFDC9;
    16'd17412: out <= 16'hFBB8;    16'd17413: out <= 16'h0058;    16'd17414: out <= 16'h03B2;    16'd17415: out <= 16'hFB4F;
    16'd17416: out <= 16'h02F3;    16'd17417: out <= 16'h02A2;    16'd17418: out <= 16'h00F0;    16'd17419: out <= 16'hFF0C;
    16'd17420: out <= 16'h032C;    16'd17421: out <= 16'hFF39;    16'd17422: out <= 16'hFF6C;    16'd17423: out <= 16'hFC52;
    16'd17424: out <= 16'hFFC5;    16'd17425: out <= 16'hFEBF;    16'd17426: out <= 16'h009A;    16'd17427: out <= 16'hFACC;
    16'd17428: out <= 16'hF8D7;    16'd17429: out <= 16'h0030;    16'd17430: out <= 16'hF88C;    16'd17431: out <= 16'h0A3F;
    16'd17432: out <= 16'h02B9;    16'd17433: out <= 16'h058A;    16'd17434: out <= 16'hF93B;    16'd17435: out <= 16'h0125;
    16'd17436: out <= 16'h088E;    16'd17437: out <= 16'hFB2D;    16'd17438: out <= 16'hFBDA;    16'd17439: out <= 16'h0414;
    16'd17440: out <= 16'h03A0;    16'd17441: out <= 16'h030B;    16'd17442: out <= 16'h00A8;    16'd17443: out <= 16'h038E;
    16'd17444: out <= 16'h0A2E;    16'd17445: out <= 16'h01A6;    16'd17446: out <= 16'h0030;    16'd17447: out <= 16'h0333;
    16'd17448: out <= 16'h0090;    16'd17449: out <= 16'h03E9;    16'd17450: out <= 16'h018B;    16'd17451: out <= 16'h076D;
    16'd17452: out <= 16'h054C;    16'd17453: out <= 16'h05AD;    16'd17454: out <= 16'h037A;    16'd17455: out <= 16'h0580;
    16'd17456: out <= 16'h0A05;    16'd17457: out <= 16'hFF2C;    16'd17458: out <= 16'h00C0;    16'd17459: out <= 16'hFFF2;
    16'd17460: out <= 16'hFDA1;    16'd17461: out <= 16'h05A3;    16'd17462: out <= 16'h08BD;    16'd17463: out <= 16'h03C2;
    16'd17464: out <= 16'h03DA;    16'd17465: out <= 16'h0104;    16'd17466: out <= 16'hFCE6;    16'd17467: out <= 16'h01B6;
    16'd17468: out <= 16'h0278;    16'd17469: out <= 16'h007A;    16'd17470: out <= 16'h0118;    16'd17471: out <= 16'h03CD;
    16'd17472: out <= 16'h043B;    16'd17473: out <= 16'h04E5;    16'd17474: out <= 16'h0420;    16'd17475: out <= 16'h024F;
    16'd17476: out <= 16'h0228;    16'd17477: out <= 16'h0231;    16'd17478: out <= 16'h04DD;    16'd17479: out <= 16'h07F2;
    16'd17480: out <= 16'hFF96;    16'd17481: out <= 16'h04CE;    16'd17482: out <= 16'hFFCB;    16'd17483: out <= 16'h04A4;
    16'd17484: out <= 16'h01A2;    16'd17485: out <= 16'h0A03;    16'd17486: out <= 16'hFDCC;    16'd17487: out <= 16'h057E;
    16'd17488: out <= 16'h0AD0;    16'd17489: out <= 16'h0396;    16'd17490: out <= 16'h0B33;    16'd17491: out <= 16'h0214;
    16'd17492: out <= 16'h08DC;    16'd17493: out <= 16'h0271;    16'd17494: out <= 16'h06BC;    16'd17495: out <= 16'h03DA;
    16'd17496: out <= 16'h0553;    16'd17497: out <= 16'h037C;    16'd17498: out <= 16'h04BD;    16'd17499: out <= 16'hFE27;
    16'd17500: out <= 16'h08BF;    16'd17501: out <= 16'h09E6;    16'd17502: out <= 16'h00EE;    16'd17503: out <= 16'hFD75;
    16'd17504: out <= 16'h01AC;    16'd17505: out <= 16'h016B;    16'd17506: out <= 16'h040D;    16'd17507: out <= 16'h030D;
    16'd17508: out <= 16'h04F8;    16'd17509: out <= 16'h0801;    16'd17510: out <= 16'h099F;    16'd17511: out <= 16'h02E6;
    16'd17512: out <= 16'h056C;    16'd17513: out <= 16'h059B;    16'd17514: out <= 16'hFCEC;    16'd17515: out <= 16'h003E;
    16'd17516: out <= 16'h04ED;    16'd17517: out <= 16'h05C3;    16'd17518: out <= 16'hFFED;    16'd17519: out <= 16'h053E;
    16'd17520: out <= 16'h0664;    16'd17521: out <= 16'h00F1;    16'd17522: out <= 16'h0683;    16'd17523: out <= 16'h0352;
    16'd17524: out <= 16'h0500;    16'd17525: out <= 16'h00DC;    16'd17526: out <= 16'h0D31;    16'd17527: out <= 16'h056E;
    16'd17528: out <= 16'hFE70;    16'd17529: out <= 16'h0828;    16'd17530: out <= 16'hFF88;    16'd17531: out <= 16'h0683;
    16'd17532: out <= 16'h0820;    16'd17533: out <= 16'hFED2;    16'd17534: out <= 16'h08D4;    16'd17535: out <= 16'h03DA;
    16'd17536: out <= 16'h035E;    16'd17537: out <= 16'h0570;    16'd17538: out <= 16'h0701;    16'd17539: out <= 16'h031D;
    16'd17540: out <= 16'h0147;    16'd17541: out <= 16'h07E6;    16'd17542: out <= 16'h00B3;    16'd17543: out <= 16'h0796;
    16'd17544: out <= 16'h0259;    16'd17545: out <= 16'h06A9;    16'd17546: out <= 16'h03FA;    16'd17547: out <= 16'h0331;
    16'd17548: out <= 16'h0499;    16'd17549: out <= 16'h05D3;    16'd17550: out <= 16'hFF98;    16'd17551: out <= 16'h056F;
    16'd17552: out <= 16'h0008;    16'd17553: out <= 16'h067A;    16'd17554: out <= 16'h0181;    16'd17555: out <= 16'h0646;
    16'd17556: out <= 16'h0626;    16'd17557: out <= 16'h04E4;    16'd17558: out <= 16'h0321;    16'd17559: out <= 16'h0A9C;
    16'd17560: out <= 16'h031E;    16'd17561: out <= 16'h010D;    16'd17562: out <= 16'h0722;    16'd17563: out <= 16'h01B5;
    16'd17564: out <= 16'h0856;    16'd17565: out <= 16'h0A0A;    16'd17566: out <= 16'h06F1;    16'd17567: out <= 16'h0502;
    16'd17568: out <= 16'h0CDD;    16'd17569: out <= 16'h047E;    16'd17570: out <= 16'h0178;    16'd17571: out <= 16'h0946;
    16'd17572: out <= 16'h04DC;    16'd17573: out <= 16'h01DE;    16'd17574: out <= 16'hFFDB;    16'd17575: out <= 16'h0622;
    16'd17576: out <= 16'h0445;    16'd17577: out <= 16'h0410;    16'd17578: out <= 16'hFB59;    16'd17579: out <= 16'hFEE0;
    16'd17580: out <= 16'h04B9;    16'd17581: out <= 16'h07DC;    16'd17582: out <= 16'h0310;    16'd17583: out <= 16'h096F;
    16'd17584: out <= 16'h0671;    16'd17585: out <= 16'h077B;    16'd17586: out <= 16'h069C;    16'd17587: out <= 16'h02DC;
    16'd17588: out <= 16'h0004;    16'd17589: out <= 16'h096F;    16'd17590: out <= 16'h0026;    16'd17591: out <= 16'h04CE;
    16'd17592: out <= 16'h04A4;    16'd17593: out <= 16'h0743;    16'd17594: out <= 16'h0009;    16'd17595: out <= 16'h001F;
    16'd17596: out <= 16'h0888;    16'd17597: out <= 16'h022F;    16'd17598: out <= 16'h03A5;    16'd17599: out <= 16'h046C;
    16'd17600: out <= 16'h0370;    16'd17601: out <= 16'h06BE;    16'd17602: out <= 16'h0723;    16'd17603: out <= 16'h0175;
    16'd17604: out <= 16'h0503;    16'd17605: out <= 16'hFF39;    16'd17606: out <= 16'h02CF;    16'd17607: out <= 16'h0499;
    16'd17608: out <= 16'h0359;    16'd17609: out <= 16'h0C03;    16'd17610: out <= 16'h0410;    16'd17611: out <= 16'h0612;
    16'd17612: out <= 16'h08C5;    16'd17613: out <= 16'hFFA7;    16'd17614: out <= 16'h0711;    16'd17615: out <= 16'hFBB2;
    16'd17616: out <= 16'h04A6;    16'd17617: out <= 16'h0264;    16'd17618: out <= 16'h0725;    16'd17619: out <= 16'h09C8;
    16'd17620: out <= 16'hFE10;    16'd17621: out <= 16'h0222;    16'd17622: out <= 16'h04A1;    16'd17623: out <= 16'h01FD;
    16'd17624: out <= 16'h0833;    16'd17625: out <= 16'h0157;    16'd17626: out <= 16'h05CD;    16'd17627: out <= 16'hFE49;
    16'd17628: out <= 16'hF8F0;    16'd17629: out <= 16'hF2D8;    16'd17630: out <= 16'h0704;    16'd17631: out <= 16'h0366;
    16'd17632: out <= 16'h00DD;    16'd17633: out <= 16'hFECF;    16'd17634: out <= 16'hFECB;    16'd17635: out <= 16'h00B5;
    16'd17636: out <= 16'hFE07;    16'd17637: out <= 16'h03F8;    16'd17638: out <= 16'h00AD;    16'd17639: out <= 16'hF94F;
    16'd17640: out <= 16'hFD12;    16'd17641: out <= 16'h0488;    16'd17642: out <= 16'hFACC;    16'd17643: out <= 16'h0780;
    16'd17644: out <= 16'hFF85;    16'd17645: out <= 16'h009A;    16'd17646: out <= 16'h0375;    16'd17647: out <= 16'hF68D;
    16'd17648: out <= 16'h040A;    16'd17649: out <= 16'h0261;    16'd17650: out <= 16'h0102;    16'd17651: out <= 16'h06F9;
    16'd17652: out <= 16'hFEDB;    16'd17653: out <= 16'hFFE6;    16'd17654: out <= 16'hFD97;    16'd17655: out <= 16'h0727;
    16'd17656: out <= 16'hFFF0;    16'd17657: out <= 16'h04CC;    16'd17658: out <= 16'h013A;    16'd17659: out <= 16'h030D;
    16'd17660: out <= 16'h00F1;    16'd17661: out <= 16'hF836;    16'd17662: out <= 16'hFF2E;    16'd17663: out <= 16'h0237;
    16'd17664: out <= 16'h0169;    16'd17665: out <= 16'h01AC;    16'd17666: out <= 16'h01FB;    16'd17667: out <= 16'hFE19;
    16'd17668: out <= 16'hFFAE;    16'd17669: out <= 16'hFCCA;    16'd17670: out <= 16'hFCD4;    16'd17671: out <= 16'hF6CD;
    16'd17672: out <= 16'h03B9;    16'd17673: out <= 16'hFD1B;    16'd17674: out <= 16'hFFDA;    16'd17675: out <= 16'h024D;
    16'd17676: out <= 16'hF6CA;    16'd17677: out <= 16'h032F;    16'd17678: out <= 16'h067B;    16'd17679: out <= 16'h0243;
    16'd17680: out <= 16'h052B;    16'd17681: out <= 16'hFE4A;    16'd17682: out <= 16'hFAE6;    16'd17683: out <= 16'hFECE;
    16'd17684: out <= 16'hFA3A;    16'd17685: out <= 16'h0453;    16'd17686: out <= 16'h0150;    16'd17687: out <= 16'hFB9C;
    16'd17688: out <= 16'h024D;    16'd17689: out <= 16'h0358;    16'd17690: out <= 16'hFFEA;    16'd17691: out <= 16'hFB44;
    16'd17692: out <= 16'h0741;    16'd17693: out <= 16'h05DB;    16'd17694: out <= 16'h0301;    16'd17695: out <= 16'h0675;
    16'd17696: out <= 16'h064E;    16'd17697: out <= 16'h0556;    16'd17698: out <= 16'h01A9;    16'd17699: out <= 16'h06D6;
    16'd17700: out <= 16'h0082;    16'd17701: out <= 16'hFAB1;    16'd17702: out <= 16'h01B0;    16'd17703: out <= 16'h029D;
    16'd17704: out <= 16'h00EA;    16'd17705: out <= 16'h0BD6;    16'd17706: out <= 16'h09A9;    16'd17707: out <= 16'h0521;
    16'd17708: out <= 16'h093E;    16'd17709: out <= 16'h0498;    16'd17710: out <= 16'hFDD1;    16'd17711: out <= 16'hFCEC;
    16'd17712: out <= 16'hFE3F;    16'd17713: out <= 16'h09A6;    16'd17714: out <= 16'h03D6;    16'd17715: out <= 16'h0016;
    16'd17716: out <= 16'h0197;    16'd17717: out <= 16'h0438;    16'd17718: out <= 16'h02C1;    16'd17719: out <= 16'h0ADA;
    16'd17720: out <= 16'h0451;    16'd17721: out <= 16'h000C;    16'd17722: out <= 16'h08A9;    16'd17723: out <= 16'h077A;
    16'd17724: out <= 16'h0205;    16'd17725: out <= 16'h00EC;    16'd17726: out <= 16'h03A6;    16'd17727: out <= 16'h0161;
    16'd17728: out <= 16'h05C5;    16'd17729: out <= 16'h071B;    16'd17730: out <= 16'h040A;    16'd17731: out <= 16'h076F;
    16'd17732: out <= 16'h08C4;    16'd17733: out <= 16'h076C;    16'd17734: out <= 16'h0425;    16'd17735: out <= 16'h077B;
    16'd17736: out <= 16'h0210;    16'd17737: out <= 16'h0345;    16'd17738: out <= 16'h05D7;    16'd17739: out <= 16'h00AC;
    16'd17740: out <= 16'h0286;    16'd17741: out <= 16'hFE48;    16'd17742: out <= 16'h009E;    16'd17743: out <= 16'h097B;
    16'd17744: out <= 16'h05DD;    16'd17745: out <= 16'h00A5;    16'd17746: out <= 16'h0576;    16'd17747: out <= 16'h0035;
    16'd17748: out <= 16'h0893;    16'd17749: out <= 16'h0667;    16'd17750: out <= 16'hFCC0;    16'd17751: out <= 16'hFC54;
    16'd17752: out <= 16'hFDCB;    16'd17753: out <= 16'h092D;    16'd17754: out <= 16'h08D9;    16'd17755: out <= 16'h0447;
    16'd17756: out <= 16'h0828;    16'd17757: out <= 16'h06FE;    16'd17758: out <= 16'h0648;    16'd17759: out <= 16'h05CA;
    16'd17760: out <= 16'h0173;    16'd17761: out <= 16'h065A;    16'd17762: out <= 16'h0976;    16'd17763: out <= 16'h0463;
    16'd17764: out <= 16'h04B2;    16'd17765: out <= 16'h063E;    16'd17766: out <= 16'h0845;    16'd17767: out <= 16'h068D;
    16'd17768: out <= 16'h0731;    16'd17769: out <= 16'h0033;    16'd17770: out <= 16'h02F7;    16'd17771: out <= 16'h06ED;
    16'd17772: out <= 16'h04F3;    16'd17773: out <= 16'h0535;    16'd17774: out <= 16'h03F8;    16'd17775: out <= 16'h08C3;
    16'd17776: out <= 16'h0504;    16'd17777: out <= 16'h05BF;    16'd17778: out <= 16'h035F;    16'd17779: out <= 16'hFE7B;
    16'd17780: out <= 16'h0CF3;    16'd17781: out <= 16'h067A;    16'd17782: out <= 16'h059E;    16'd17783: out <= 16'hFCDA;
    16'd17784: out <= 16'h0545;    16'd17785: out <= 16'h0084;    16'd17786: out <= 16'h00C3;    16'd17787: out <= 16'h02D8;
    16'd17788: out <= 16'hFEC1;    16'd17789: out <= 16'h0414;    16'd17790: out <= 16'h026E;    16'd17791: out <= 16'h0642;
    16'd17792: out <= 16'h0A87;    16'd17793: out <= 16'h0485;    16'd17794: out <= 16'h06B4;    16'd17795: out <= 16'h017E;
    16'd17796: out <= 16'h0D3B;    16'd17797: out <= 16'h05DB;    16'd17798: out <= 16'h04A4;    16'd17799: out <= 16'h037D;
    16'd17800: out <= 16'h04CF;    16'd17801: out <= 16'h0734;    16'd17802: out <= 16'h054A;    16'd17803: out <= 16'hFDE2;
    16'd17804: out <= 16'h0289;    16'd17805: out <= 16'hFD1C;    16'd17806: out <= 16'h0492;    16'd17807: out <= 16'h0832;
    16'd17808: out <= 16'h02EE;    16'd17809: out <= 16'h05E4;    16'd17810: out <= 16'h0689;    16'd17811: out <= 16'h039B;
    16'd17812: out <= 16'h0B5B;    16'd17813: out <= 16'h054C;    16'd17814: out <= 16'h0080;    16'd17815: out <= 16'h0677;
    16'd17816: out <= 16'h0643;    16'd17817: out <= 16'h0486;    16'd17818: out <= 16'hFD83;    16'd17819: out <= 16'h0A6A;
    16'd17820: out <= 16'h0583;    16'd17821: out <= 16'h02DF;    16'd17822: out <= 16'h06C9;    16'd17823: out <= 16'hFF03;
    16'd17824: out <= 16'hFF0E;    16'd17825: out <= 16'hFE01;    16'd17826: out <= 16'h02BE;    16'd17827: out <= 16'h0597;
    16'd17828: out <= 16'h0157;    16'd17829: out <= 16'h03CA;    16'd17830: out <= 16'h010B;    16'd17831: out <= 16'h0586;
    16'd17832: out <= 16'h0502;    16'd17833: out <= 16'h0523;    16'd17834: out <= 16'h07DE;    16'd17835: out <= 16'hFC5C;
    16'd17836: out <= 16'h070C;    16'd17837: out <= 16'h04D7;    16'd17838: out <= 16'hFB7F;    16'd17839: out <= 16'h0769;
    16'd17840: out <= 16'h0449;    16'd17841: out <= 16'h0069;    16'd17842: out <= 16'h0674;    16'd17843: out <= 16'h018B;
    16'd17844: out <= 16'h061C;    16'd17845: out <= 16'h02FE;    16'd17846: out <= 16'h0358;    16'd17847: out <= 16'h04CB;
    16'd17848: out <= 16'h06AD;    16'd17849: out <= 16'hFFDF;    16'd17850: out <= 16'h05E8;    16'd17851: out <= 16'h004D;
    16'd17852: out <= 16'hFF60;    16'd17853: out <= 16'h01BF;    16'd17854: out <= 16'h0209;    16'd17855: out <= 16'h0721;
    16'd17856: out <= 16'h00DF;    16'd17857: out <= 16'hFF7F;    16'd17858: out <= 16'hFF0B;    16'd17859: out <= 16'h0352;
    16'd17860: out <= 16'h0584;    16'd17861: out <= 16'h0580;    16'd17862: out <= 16'hFF6F;    16'd17863: out <= 16'h02A2;
    16'd17864: out <= 16'h0A30;    16'd17865: out <= 16'h07AB;    16'd17866: out <= 16'h02A1;    16'd17867: out <= 16'h082C;
    16'd17868: out <= 16'h0357;    16'd17869: out <= 16'hFB2E;    16'd17870: out <= 16'h0441;    16'd17871: out <= 16'h03E7;
    16'd17872: out <= 16'hFF4D;    16'd17873: out <= 16'h05F1;    16'd17874: out <= 16'hFBD5;    16'd17875: out <= 16'h0818;
    16'd17876: out <= 16'h0268;    16'd17877: out <= 16'h011C;    16'd17878: out <= 16'hFF9E;    16'd17879: out <= 16'h0189;
    16'd17880: out <= 16'h0254;    16'd17881: out <= 16'hFFF5;    16'd17882: out <= 16'h0158;    16'd17883: out <= 16'hFED2;
    16'd17884: out <= 16'h0239;    16'd17885: out <= 16'h0374;    16'd17886: out <= 16'hF62C;    16'd17887: out <= 16'h02FC;
    16'd17888: out <= 16'h0754;    16'd17889: out <= 16'hFDB5;    16'd17890: out <= 16'hFFE6;    16'd17891: out <= 16'h02AD;
    16'd17892: out <= 16'h0080;    16'd17893: out <= 16'hFDB8;    16'd17894: out <= 16'h0028;    16'd17895: out <= 16'h00E7;
    16'd17896: out <= 16'hFB61;    16'd17897: out <= 16'hFEFB;    16'd17898: out <= 16'hFE1A;    16'd17899: out <= 16'hFF55;
    16'd17900: out <= 16'hF9EE;    16'd17901: out <= 16'h01C7;    16'd17902: out <= 16'h031E;    16'd17903: out <= 16'h05B8;
    16'd17904: out <= 16'h024D;    16'd17905: out <= 16'hFC22;    16'd17906: out <= 16'h004D;    16'd17907: out <= 16'h030B;
    16'd17908: out <= 16'h00AD;    16'd17909: out <= 16'hFF7B;    16'd17910: out <= 16'h04C6;    16'd17911: out <= 16'hFF61;
    16'd17912: out <= 16'hFD60;    16'd17913: out <= 16'hFE4A;    16'd17914: out <= 16'h06BC;    16'd17915: out <= 16'h0530;
    16'd17916: out <= 16'hFD83;    16'd17917: out <= 16'h0138;    16'd17918: out <= 16'h0102;    16'd17919: out <= 16'hFF0F;
    16'd17920: out <= 16'h038C;    16'd17921: out <= 16'hFF4E;    16'd17922: out <= 16'h080B;    16'd17923: out <= 16'h0365;
    16'd17924: out <= 16'h019C;    16'd17925: out <= 16'hFA9B;    16'd17926: out <= 16'h045B;    16'd17927: out <= 16'hFF1F;
    16'd17928: out <= 16'hFE96;    16'd17929: out <= 16'h03E6;    16'd17930: out <= 16'hFF28;    16'd17931: out <= 16'hFF8E;
    16'd17932: out <= 16'hFB30;    16'd17933: out <= 16'hFDA7;    16'd17934: out <= 16'hFBCD;    16'd17935: out <= 16'hFFC1;
    16'd17936: out <= 16'h0171;    16'd17937: out <= 16'hFC2A;    16'd17938: out <= 16'h0083;    16'd17939: out <= 16'h00D0;
    16'd17940: out <= 16'h0331;    16'd17941: out <= 16'hFC68;    16'd17942: out <= 16'h0153;    16'd17943: out <= 16'hFDF4;
    16'd17944: out <= 16'h04B0;    16'd17945: out <= 16'hFFD4;    16'd17946: out <= 16'hFF8B;    16'd17947: out <= 16'hFDBC;
    16'd17948: out <= 16'h034C;    16'd17949: out <= 16'h09F6;    16'd17950: out <= 16'h0285;    16'd17951: out <= 16'hFBF3;
    16'd17952: out <= 16'h047A;    16'd17953: out <= 16'h00B9;    16'd17954: out <= 16'h0724;    16'd17955: out <= 16'h010D;
    16'd17956: out <= 16'h031C;    16'd17957: out <= 16'h0168;    16'd17958: out <= 16'h000F;    16'd17959: out <= 16'h00F3;
    16'd17960: out <= 16'h036E;    16'd17961: out <= 16'h058D;    16'd17962: out <= 16'h0881;    16'd17963: out <= 16'hFD6A;
    16'd17964: out <= 16'h091D;    16'd17965: out <= 16'hFCB8;    16'd17966: out <= 16'h0477;    16'd17967: out <= 16'h00BC;
    16'd17968: out <= 16'h05CA;    16'd17969: out <= 16'h0660;    16'd17970: out <= 16'h03FF;    16'd17971: out <= 16'h0855;
    16'd17972: out <= 16'h01D8;    16'd17973: out <= 16'h0264;    16'd17974: out <= 16'hFE69;    16'd17975: out <= 16'h0546;
    16'd17976: out <= 16'h05D6;    16'd17977: out <= 16'h00DB;    16'd17978: out <= 16'h02E1;    16'd17979: out <= 16'h0AB6;
    16'd17980: out <= 16'hFE35;    16'd17981: out <= 16'hFF36;    16'd17982: out <= 16'h06E1;    16'd17983: out <= 16'h0002;
    16'd17984: out <= 16'h0233;    16'd17985: out <= 16'h05BA;    16'd17986: out <= 16'hFE70;    16'd17987: out <= 16'hFFA9;
    16'd17988: out <= 16'h0781;    16'd17989: out <= 16'h0071;    16'd17990: out <= 16'h0362;    16'd17991: out <= 16'h0A4F;
    16'd17992: out <= 16'h0470;    16'd17993: out <= 16'hFF4C;    16'd17994: out <= 16'h077A;    16'd17995: out <= 16'h01ED;
    16'd17996: out <= 16'h011A;    16'd17997: out <= 16'h04DC;    16'd17998: out <= 16'h011A;    16'd17999: out <= 16'h00D8;
    16'd18000: out <= 16'h05FB;    16'd18001: out <= 16'hFBA5;    16'd18002: out <= 16'h02C4;    16'd18003: out <= 16'hFE25;
    16'd18004: out <= 16'h08D4;    16'd18005: out <= 16'h00D4;    16'd18006: out <= 16'hFF4E;    16'd18007: out <= 16'h03ED;
    16'd18008: out <= 16'h0591;    16'd18009: out <= 16'h07AA;    16'd18010: out <= 16'h071D;    16'd18011: out <= 16'h02AF;
    16'd18012: out <= 16'h00D3;    16'd18013: out <= 16'hFED3;    16'd18014: out <= 16'h04A1;    16'd18015: out <= 16'h0239;
    16'd18016: out <= 16'h0681;    16'd18017: out <= 16'h015A;    16'd18018: out <= 16'hFB6A;    16'd18019: out <= 16'h0340;
    16'd18020: out <= 16'hFF8D;    16'd18021: out <= 16'h06EB;    16'd18022: out <= 16'h087B;    16'd18023: out <= 16'h0637;
    16'd18024: out <= 16'hFEF5;    16'd18025: out <= 16'h0BE2;    16'd18026: out <= 16'h023D;    16'd18027: out <= 16'h0C09;
    16'd18028: out <= 16'h11C9;    16'd18029: out <= 16'h0A59;    16'd18030: out <= 16'h025E;    16'd18031: out <= 16'h0297;
    16'd18032: out <= 16'h0970;    16'd18033: out <= 16'h0197;    16'd18034: out <= 16'h0714;    16'd18035: out <= 16'hFE1B;
    16'd18036: out <= 16'h040C;    16'd18037: out <= 16'h0432;    16'd18038: out <= 16'h0317;    16'd18039: out <= 16'h058C;
    16'd18040: out <= 16'h033C;    16'd18041: out <= 16'h06FB;    16'd18042: out <= 16'h083C;    16'd18043: out <= 16'h0489;
    16'd18044: out <= 16'h050A;    16'd18045: out <= 16'hFD1E;    16'd18046: out <= 16'h0465;    16'd18047: out <= 16'h083C;
    16'd18048: out <= 16'h02D5;    16'd18049: out <= 16'hFDB9;    16'd18050: out <= 16'h0252;    16'd18051: out <= 16'h0154;
    16'd18052: out <= 16'hFFEF;    16'd18053: out <= 16'h07AF;    16'd18054: out <= 16'h0320;    16'd18055: out <= 16'h01BC;
    16'd18056: out <= 16'hF92B;    16'd18057: out <= 16'h04A7;    16'd18058: out <= 16'h0925;    16'd18059: out <= 16'h0734;
    16'd18060: out <= 16'h07CD;    16'd18061: out <= 16'h01FC;    16'd18062: out <= 16'h0972;    16'd18063: out <= 16'h0732;
    16'd18064: out <= 16'h0595;    16'd18065: out <= 16'h070B;    16'd18066: out <= 16'h06B4;    16'd18067: out <= 16'hFE48;
    16'd18068: out <= 16'h0101;    16'd18069: out <= 16'h0551;    16'd18070: out <= 16'h033B;    16'd18071: out <= 16'h03A8;
    16'd18072: out <= 16'h0B3F;    16'd18073: out <= 16'h06E0;    16'd18074: out <= 16'h01AE;    16'd18075: out <= 16'h0059;
    16'd18076: out <= 16'h00B5;    16'd18077: out <= 16'h0197;    16'd18078: out <= 16'hFE6F;    16'd18079: out <= 16'h0311;
    16'd18080: out <= 16'h007A;    16'd18081: out <= 16'h0257;    16'd18082: out <= 16'h0697;    16'd18083: out <= 16'hFE0E;
    16'd18084: out <= 16'hFF52;    16'd18085: out <= 16'hFF83;    16'd18086: out <= 16'h0336;    16'd18087: out <= 16'hFE2F;
    16'd18088: out <= 16'h0656;    16'd18089: out <= 16'hFA5A;    16'd18090: out <= 16'h0444;    16'd18091: out <= 16'h0964;
    16'd18092: out <= 16'hFB74;    16'd18093: out <= 16'h04DB;    16'd18094: out <= 16'h0434;    16'd18095: out <= 16'h0258;
    16'd18096: out <= 16'h0533;    16'd18097: out <= 16'h05AF;    16'd18098: out <= 16'h06B9;    16'd18099: out <= 16'h049B;
    16'd18100: out <= 16'h01F7;    16'd18101: out <= 16'h05A1;    16'd18102: out <= 16'h0888;    16'd18103: out <= 16'h0629;
    16'd18104: out <= 16'h001A;    16'd18105: out <= 16'hFEDC;    16'd18106: out <= 16'h0A39;    16'd18107: out <= 16'h017A;
    16'd18108: out <= 16'hFFC8;    16'd18109: out <= 16'h0165;    16'd18110: out <= 16'h00EA;    16'd18111: out <= 16'h064D;
    16'd18112: out <= 16'h06E7;    16'd18113: out <= 16'h08EF;    16'd18114: out <= 16'h076C;    16'd18115: out <= 16'h0804;
    16'd18116: out <= 16'h0745;    16'd18117: out <= 16'h01DC;    16'd18118: out <= 16'h0C66;    16'd18119: out <= 16'hFB86;
    16'd18120: out <= 16'hF9D8;    16'd18121: out <= 16'hFE9B;    16'd18122: out <= 16'hF9DF;    16'd18123: out <= 16'h01B2;
    16'd18124: out <= 16'h0586;    16'd18125: out <= 16'h07A5;    16'd18126: out <= 16'h026F;    16'd18127: out <= 16'h081F;
    16'd18128: out <= 16'h065A;    16'd18129: out <= 16'h02CC;    16'd18130: out <= 16'h0E56;    16'd18131: out <= 16'h0822;
    16'd18132: out <= 16'h0386;    16'd18133: out <= 16'hFF1D;    16'd18134: out <= 16'h036B;    16'd18135: out <= 16'hFB6F;
    16'd18136: out <= 16'h0573;    16'd18137: out <= 16'h0210;    16'd18138: out <= 16'h038D;    16'd18139: out <= 16'hFF8B;
    16'd18140: out <= 16'hFCF3;    16'd18141: out <= 16'hF9E5;    16'd18142: out <= 16'h04E6;    16'd18143: out <= 16'hF77C;
    16'd18144: out <= 16'h0738;    16'd18145: out <= 16'h05B5;    16'd18146: out <= 16'h07A3;    16'd18147: out <= 16'h0071;
    16'd18148: out <= 16'hFCA0;    16'd18149: out <= 16'hFFFF;    16'd18150: out <= 16'hFEA8;    16'd18151: out <= 16'h0058;
    16'd18152: out <= 16'h03B0;    16'd18153: out <= 16'h04B5;    16'd18154: out <= 16'h093E;    16'd18155: out <= 16'h03EA;
    16'd18156: out <= 16'hFB9A;    16'd18157: out <= 16'h0318;    16'd18158: out <= 16'hF9A2;    16'd18159: out <= 16'hFB16;
    16'd18160: out <= 16'h03C7;    16'd18161: out <= 16'h0058;    16'd18162: out <= 16'h011E;    16'd18163: out <= 16'hF84F;
    16'd18164: out <= 16'hFB89;    16'd18165: out <= 16'h0029;    16'd18166: out <= 16'h06BE;    16'd18167: out <= 16'h0371;
    16'd18168: out <= 16'hFF32;    16'd18169: out <= 16'h040C;    16'd18170: out <= 16'hFA3D;    16'd18171: out <= 16'hFF93;
    16'd18172: out <= 16'hFD42;    16'd18173: out <= 16'h0252;    16'd18174: out <= 16'h07E5;    16'd18175: out <= 16'hFCF8;
    16'd18176: out <= 16'h0353;    16'd18177: out <= 16'hF84A;    16'd18178: out <= 16'hFA8C;    16'd18179: out <= 16'h0618;
    16'd18180: out <= 16'h025D;    16'd18181: out <= 16'hFD73;    16'd18182: out <= 16'hFC2B;    16'd18183: out <= 16'h01E2;
    16'd18184: out <= 16'h0148;    16'd18185: out <= 16'hFA9D;    16'd18186: out <= 16'hFE8E;    16'd18187: out <= 16'h01A9;
    16'd18188: out <= 16'hFE53;    16'd18189: out <= 16'h00F6;    16'd18190: out <= 16'h03EB;    16'd18191: out <= 16'hFEAC;
    16'd18192: out <= 16'h01BE;    16'd18193: out <= 16'hF9E6;    16'd18194: out <= 16'h02B3;    16'd18195: out <= 16'hFCAE;
    16'd18196: out <= 16'hFF58;    16'd18197: out <= 16'hFCBB;    16'd18198: out <= 16'hFD35;    16'd18199: out <= 16'h01C8;
    16'd18200: out <= 16'h03F2;    16'd18201: out <= 16'hFEEE;    16'd18202: out <= 16'h078B;    16'd18203: out <= 16'h010B;
    16'd18204: out <= 16'h0284;    16'd18205: out <= 16'h067E;    16'd18206: out <= 16'h0018;    16'd18207: out <= 16'hFEF5;
    16'd18208: out <= 16'h04D3;    16'd18209: out <= 16'h002D;    16'd18210: out <= 16'h0657;    16'd18211: out <= 16'h04DC;
    16'd18212: out <= 16'h027F;    16'd18213: out <= 16'h0473;    16'd18214: out <= 16'h0920;    16'd18215: out <= 16'h0266;
    16'd18216: out <= 16'h0371;    16'd18217: out <= 16'hFDE7;    16'd18218: out <= 16'h04B3;    16'd18219: out <= 16'h09C2;
    16'd18220: out <= 16'h0997;    16'd18221: out <= 16'h06DD;    16'd18222: out <= 16'h018B;    16'd18223: out <= 16'h052C;
    16'd18224: out <= 16'h0346;    16'd18225: out <= 16'h0A4A;    16'd18226: out <= 16'hFF53;    16'd18227: out <= 16'hFD2F;
    16'd18228: out <= 16'h04D5;    16'd18229: out <= 16'h0319;    16'd18230: out <= 16'h0C18;    16'd18231: out <= 16'h0305;
    16'd18232: out <= 16'h0639;    16'd18233: out <= 16'h038E;    16'd18234: out <= 16'h0523;    16'd18235: out <= 16'h012F;
    16'd18236: out <= 16'h0044;    16'd18237: out <= 16'h047C;    16'd18238: out <= 16'h021C;    16'd18239: out <= 16'h02DF;
    16'd18240: out <= 16'h047F;    16'd18241: out <= 16'h02D6;    16'd18242: out <= 16'hFF18;    16'd18243: out <= 16'h0880;
    16'd18244: out <= 16'h0776;    16'd18245: out <= 16'h00DC;    16'd18246: out <= 16'h057B;    16'd18247: out <= 16'h038F;
    16'd18248: out <= 16'hFFA5;    16'd18249: out <= 16'h03C2;    16'd18250: out <= 16'h0882;    16'd18251: out <= 16'h056F;
    16'd18252: out <= 16'hFFFF;    16'd18253: out <= 16'h0B0F;    16'd18254: out <= 16'h0243;    16'd18255: out <= 16'hFDF7;
    16'd18256: out <= 16'h0142;    16'd18257: out <= 16'h02D0;    16'd18258: out <= 16'hFD39;    16'd18259: out <= 16'h0608;
    16'd18260: out <= 16'h040A;    16'd18261: out <= 16'hFE14;    16'd18262: out <= 16'hFF4C;    16'd18263: out <= 16'h0042;
    16'd18264: out <= 16'h0763;    16'd18265: out <= 16'h0990;    16'd18266: out <= 16'h08EF;    16'd18267: out <= 16'h04D1;
    16'd18268: out <= 16'hFF2B;    16'd18269: out <= 16'h043C;    16'd18270: out <= 16'h035E;    16'd18271: out <= 16'h0309;
    16'd18272: out <= 16'h07DC;    16'd18273: out <= 16'h0502;    16'd18274: out <= 16'h0253;    16'd18275: out <= 16'h02CE;
    16'd18276: out <= 16'h0219;    16'd18277: out <= 16'hFF70;    16'd18278: out <= 16'h045E;    16'd18279: out <= 16'h01F7;
    16'd18280: out <= 16'h0159;    16'd18281: out <= 16'h03C7;    16'd18282: out <= 16'h08BF;    16'd18283: out <= 16'h02D1;
    16'd18284: out <= 16'h080C;    16'd18285: out <= 16'h083D;    16'd18286: out <= 16'h08CD;    16'd18287: out <= 16'h07E1;
    16'd18288: out <= 16'hFDD6;    16'd18289: out <= 16'hFFEE;    16'd18290: out <= 16'h00BF;    16'd18291: out <= 16'h02DC;
    16'd18292: out <= 16'h055A;    16'd18293: out <= 16'hFF2F;    16'd18294: out <= 16'h0874;    16'd18295: out <= 16'h0058;
    16'd18296: out <= 16'h090E;    16'd18297: out <= 16'h03AE;    16'd18298: out <= 16'h0139;    16'd18299: out <= 16'hFACC;
    16'd18300: out <= 16'hFF5E;    16'd18301: out <= 16'h0456;    16'd18302: out <= 16'h070D;    16'd18303: out <= 16'hFFC9;
    16'd18304: out <= 16'h06B6;    16'd18305: out <= 16'h0307;    16'd18306: out <= 16'hFE97;    16'd18307: out <= 16'hFFA2;
    16'd18308: out <= 16'h0096;    16'd18309: out <= 16'h0211;    16'd18310: out <= 16'h050A;    16'd18311: out <= 16'hFFF9;
    16'd18312: out <= 16'h030A;    16'd18313: out <= 16'h0D72;    16'd18314: out <= 16'h0555;    16'd18315: out <= 16'h097B;
    16'd18316: out <= 16'h053C;    16'd18317: out <= 16'h0470;    16'd18318: out <= 16'h03FF;    16'd18319: out <= 16'h05A7;
    16'd18320: out <= 16'h03CD;    16'd18321: out <= 16'h086C;    16'd18322: out <= 16'h02A8;    16'd18323: out <= 16'h06F7;
    16'd18324: out <= 16'h0ADE;    16'd18325: out <= 16'h00E9;    16'd18326: out <= 16'hFD40;    16'd18327: out <= 16'h062D;
    16'd18328: out <= 16'h0541;    16'd18329: out <= 16'h06A4;    16'd18330: out <= 16'h038D;    16'd18331: out <= 16'h04F5;
    16'd18332: out <= 16'hFE9A;    16'd18333: out <= 16'h0699;    16'd18334: out <= 16'h00EF;    16'd18335: out <= 16'h0676;
    16'd18336: out <= 16'h003B;    16'd18337: out <= 16'h0443;    16'd18338: out <= 16'h0400;    16'd18339: out <= 16'h020E;
    16'd18340: out <= 16'h06BE;    16'd18341: out <= 16'h03ED;    16'd18342: out <= 16'hFFEB;    16'd18343: out <= 16'h0471;
    16'd18344: out <= 16'h0488;    16'd18345: out <= 16'h09F9;    16'd18346: out <= 16'h0868;    16'd18347: out <= 16'h0770;
    16'd18348: out <= 16'h06DB;    16'd18349: out <= 16'h0BDE;    16'd18350: out <= 16'hFEA5;    16'd18351: out <= 16'h011B;
    16'd18352: out <= 16'hFFA9;    16'd18353: out <= 16'h0800;    16'd18354: out <= 16'h02DC;    16'd18355: out <= 16'h048A;
    16'd18356: out <= 16'h05B1;    16'd18357: out <= 16'h033E;    16'd18358: out <= 16'h02E2;    16'd18359: out <= 16'h02B6;
    16'd18360: out <= 16'h07CC;    16'd18361: out <= 16'hFDDB;    16'd18362: out <= 16'h0AD4;    16'd18363: out <= 16'h015B;
    16'd18364: out <= 16'h02F9;    16'd18365: out <= 16'h09BD;    16'd18366: out <= 16'h00F8;    16'd18367: out <= 16'h0684;
    16'd18368: out <= 16'hFD64;    16'd18369: out <= 16'h017F;    16'd18370: out <= 16'h06D3;    16'd18371: out <= 16'hFBD2;
    16'd18372: out <= 16'h0510;    16'd18373: out <= 16'h0054;    16'd18374: out <= 16'h0B80;    16'd18375: out <= 16'h044D;
    16'd18376: out <= 16'h07B0;    16'd18377: out <= 16'h02C1;    16'd18378: out <= 16'h002C;    16'd18379: out <= 16'h022F;
    16'd18380: out <= 16'h01AB;    16'd18381: out <= 16'hFDE9;    16'd18382: out <= 16'hFFDC;    16'd18383: out <= 16'h01C0;
    16'd18384: out <= 16'h02A4;    16'd18385: out <= 16'h0147;    16'd18386: out <= 16'h050A;    16'd18387: out <= 16'h0765;
    16'd18388: out <= 16'h035E;    16'd18389: out <= 16'hFEF8;    16'd18390: out <= 16'hFE7C;    16'd18391: out <= 16'h0470;
    16'd18392: out <= 16'h0596;    16'd18393: out <= 16'h0144;    16'd18394: out <= 16'h0230;    16'd18395: out <= 16'h017C;
    16'd18396: out <= 16'hFEC4;    16'd18397: out <= 16'hFDF5;    16'd18398: out <= 16'h026D;    16'd18399: out <= 16'hFB8A;
    16'd18400: out <= 16'hFEA4;    16'd18401: out <= 16'hFD35;    16'd18402: out <= 16'h0166;    16'd18403: out <= 16'h0506;
    16'd18404: out <= 16'h005C;    16'd18405: out <= 16'hFAA2;    16'd18406: out <= 16'h010F;    16'd18407: out <= 16'h02B4;
    16'd18408: out <= 16'h00D0;    16'd18409: out <= 16'hFCC0;    16'd18410: out <= 16'h01DF;    16'd18411: out <= 16'hFD22;
    16'd18412: out <= 16'h00CA;    16'd18413: out <= 16'h06AD;    16'd18414: out <= 16'hFDE9;    16'd18415: out <= 16'h03C0;
    16'd18416: out <= 16'h01FD;    16'd18417: out <= 16'hFF52;    16'd18418: out <= 16'h02EC;    16'd18419: out <= 16'hFC49;
    16'd18420: out <= 16'hFF1F;    16'd18421: out <= 16'h061A;    16'd18422: out <= 16'h0616;    16'd18423: out <= 16'hFC37;
    16'd18424: out <= 16'h01FD;    16'd18425: out <= 16'hFDF5;    16'd18426: out <= 16'hFAE5;    16'd18427: out <= 16'hF77A;
    16'd18428: out <= 16'h02EB;    16'd18429: out <= 16'hFF9C;    16'd18430: out <= 16'h02A4;    16'd18431: out <= 16'h011A;
    16'd18432: out <= 16'h0317;    16'd18433: out <= 16'hFBF5;    16'd18434: out <= 16'h00B6;    16'd18435: out <= 16'h0473;
    16'd18436: out <= 16'h0162;    16'd18437: out <= 16'h004D;    16'd18438: out <= 16'h0670;    16'd18439: out <= 16'hFDCD;
    16'd18440: out <= 16'h0388;    16'd18441: out <= 16'hFEC8;    16'd18442: out <= 16'h03C3;    16'd18443: out <= 16'hF96E;
    16'd18444: out <= 16'h0024;    16'd18445: out <= 16'hFE73;    16'd18446: out <= 16'hFF84;    16'd18447: out <= 16'hFB04;
    16'd18448: out <= 16'h05C6;    16'd18449: out <= 16'hF957;    16'd18450: out <= 16'hFF49;    16'd18451: out <= 16'h02C4;
    16'd18452: out <= 16'h0597;    16'd18453: out <= 16'h015F;    16'd18454: out <= 16'hFCDF;    16'd18455: out <= 16'hFEF4;
    16'd18456: out <= 16'hFEF3;    16'd18457: out <= 16'h019F;    16'd18458: out <= 16'hF674;    16'd18459: out <= 16'h0457;
    16'd18460: out <= 16'h0614;    16'd18461: out <= 16'h0617;    16'd18462: out <= 16'h08D0;    16'd18463: out <= 16'h0231;
    16'd18464: out <= 16'h03A4;    16'd18465: out <= 16'h01D9;    16'd18466: out <= 16'h071F;    16'd18467: out <= 16'h07CA;
    16'd18468: out <= 16'h027E;    16'd18469: out <= 16'h0646;    16'd18470: out <= 16'h067D;    16'd18471: out <= 16'h099B;
    16'd18472: out <= 16'h0910;    16'd18473: out <= 16'h024D;    16'd18474: out <= 16'h0619;    16'd18475: out <= 16'h0901;
    16'd18476: out <= 16'hFACD;    16'd18477: out <= 16'h0606;    16'd18478: out <= 16'h0A51;    16'd18479: out <= 16'h051B;
    16'd18480: out <= 16'h0645;    16'd18481: out <= 16'h040E;    16'd18482: out <= 16'h03E2;    16'd18483: out <= 16'hFFB8;
    16'd18484: out <= 16'h0315;    16'd18485: out <= 16'h0274;    16'd18486: out <= 16'h04EE;    16'd18487: out <= 16'h02E6;
    16'd18488: out <= 16'hFD47;    16'd18489: out <= 16'h03D8;    16'd18490: out <= 16'h050A;    16'd18491: out <= 16'h08E8;
    16'd18492: out <= 16'h0763;    16'd18493: out <= 16'h04EC;    16'd18494: out <= 16'h09B7;    16'd18495: out <= 16'h02E0;
    16'd18496: out <= 16'h0390;    16'd18497: out <= 16'h0586;    16'd18498: out <= 16'h044C;    16'd18499: out <= 16'h042B;
    16'd18500: out <= 16'h04C6;    16'd18501: out <= 16'hFDD6;    16'd18502: out <= 16'h0355;    16'd18503: out <= 16'h06BE;
    16'd18504: out <= 16'h0108;    16'd18505: out <= 16'h0775;    16'd18506: out <= 16'h01FB;    16'd18507: out <= 16'h0329;
    16'd18508: out <= 16'h0216;    16'd18509: out <= 16'h0678;    16'd18510: out <= 16'hFFEF;    16'd18511: out <= 16'h0412;
    16'd18512: out <= 16'h08F8;    16'd18513: out <= 16'h083A;    16'd18514: out <= 16'hFE99;    16'd18515: out <= 16'h0E6E;
    16'd18516: out <= 16'h00F1;    16'd18517: out <= 16'h06F8;    16'd18518: out <= 16'h030F;    16'd18519: out <= 16'h08F1;
    16'd18520: out <= 16'h0018;    16'd18521: out <= 16'hFBA9;    16'd18522: out <= 16'h008D;    16'd18523: out <= 16'h0541;
    16'd18524: out <= 16'h0141;    16'd18525: out <= 16'h0A2D;    16'd18526: out <= 16'h06A8;    16'd18527: out <= 16'hFFB8;
    16'd18528: out <= 16'h0958;    16'd18529: out <= 16'h08BD;    16'd18530: out <= 16'h06AB;    16'd18531: out <= 16'h02BE;
    16'd18532: out <= 16'h02FC;    16'd18533: out <= 16'h079E;    16'd18534: out <= 16'h024C;    16'd18535: out <= 16'h0830;
    16'd18536: out <= 16'h051D;    16'd18537: out <= 16'h0250;    16'd18538: out <= 16'h0489;    16'd18539: out <= 16'h0316;
    16'd18540: out <= 16'hFB7A;    16'd18541: out <= 16'hFF6B;    16'd18542: out <= 16'h0811;    16'd18543: out <= 16'h0C01;
    16'd18544: out <= 16'h0392;    16'd18545: out <= 16'h0938;    16'd18546: out <= 16'hFA7C;    16'd18547: out <= 16'h061C;
    16'd18548: out <= 16'h0127;    16'd18549: out <= 16'h0496;    16'd18550: out <= 16'h0103;    16'd18551: out <= 16'h075F;
    16'd18552: out <= 16'h097F;    16'd18553: out <= 16'h02E1;    16'd18554: out <= 16'h02AC;    16'd18555: out <= 16'hFFEA;
    16'd18556: out <= 16'hFE27;    16'd18557: out <= 16'h04CE;    16'd18558: out <= 16'h0273;    16'd18559: out <= 16'h0096;
    16'd18560: out <= 16'hFFF1;    16'd18561: out <= 16'h0138;    16'd18562: out <= 16'h0194;    16'd18563: out <= 16'h03E7;
    16'd18564: out <= 16'h027B;    16'd18565: out <= 16'h0535;    16'd18566: out <= 16'h0776;    16'd18567: out <= 16'h0349;
    16'd18568: out <= 16'hFD5F;    16'd18569: out <= 16'h067D;    16'd18570: out <= 16'h0297;    16'd18571: out <= 16'h0073;
    16'd18572: out <= 16'h0C79;    16'd18573: out <= 16'hFFA2;    16'd18574: out <= 16'h0174;    16'd18575: out <= 16'h0488;
    16'd18576: out <= 16'h076D;    16'd18577: out <= 16'h0729;    16'd18578: out <= 16'h0A5D;    16'd18579: out <= 16'h0759;
    16'd18580: out <= 16'h0730;    16'd18581: out <= 16'h01D0;    16'd18582: out <= 16'h071B;    16'd18583: out <= 16'h0627;
    16'd18584: out <= 16'h0856;    16'd18585: out <= 16'h0715;    16'd18586: out <= 16'h033B;    16'd18587: out <= 16'h02AA;
    16'd18588: out <= 16'hFCE5;    16'd18589: out <= 16'hFCA6;    16'd18590: out <= 16'h099E;    16'd18591: out <= 16'h0ADF;
    16'd18592: out <= 16'h0802;    16'd18593: out <= 16'h0B2F;    16'd18594: out <= 16'h05C0;    16'd18595: out <= 16'h0399;
    16'd18596: out <= 16'hFB1A;    16'd18597: out <= 16'hF878;    16'd18598: out <= 16'hFFF4;    16'd18599: out <= 16'h0828;
    16'd18600: out <= 16'h05D4;    16'd18601: out <= 16'h057B;    16'd18602: out <= 16'h0474;    16'd18603: out <= 16'hFFF8;
    16'd18604: out <= 16'hFF68;    16'd18605: out <= 16'h075B;    16'd18606: out <= 16'h01D3;    16'd18607: out <= 16'h0749;
    16'd18608: out <= 16'h0090;    16'd18609: out <= 16'h097A;    16'd18610: out <= 16'h06F8;    16'd18611: out <= 16'h0789;
    16'd18612: out <= 16'h082F;    16'd18613: out <= 16'h03F0;    16'd18614: out <= 16'h0124;    16'd18615: out <= 16'h065E;
    16'd18616: out <= 16'hFFAD;    16'd18617: out <= 16'h03D4;    16'd18618: out <= 16'h06C6;    16'd18619: out <= 16'h0736;
    16'd18620: out <= 16'h03AA;    16'd18621: out <= 16'h084E;    16'd18622: out <= 16'h069E;    16'd18623: out <= 16'h06EC;
    16'd18624: out <= 16'h0626;    16'd18625: out <= 16'h0323;    16'd18626: out <= 16'h054B;    16'd18627: out <= 16'h009F;
    16'd18628: out <= 16'h075C;    16'd18629: out <= 16'h01CB;    16'd18630: out <= 16'h00B6;    16'd18631: out <= 16'h09D0;
    16'd18632: out <= 16'h0428;    16'd18633: out <= 16'h04CC;    16'd18634: out <= 16'h038C;    16'd18635: out <= 16'h06D3;
    16'd18636: out <= 16'h0741;    16'd18637: out <= 16'h0C7A;    16'd18638: out <= 16'h0190;    16'd18639: out <= 16'h0021;
    16'd18640: out <= 16'h0A10;    16'd18641: out <= 16'h0942;    16'd18642: out <= 16'h02C3;    16'd18643: out <= 16'hFEC0;
    16'd18644: out <= 16'h0454;    16'd18645: out <= 16'h087F;    16'd18646: out <= 16'h04C3;    16'd18647: out <= 16'h0A7A;
    16'd18648: out <= 16'h050A;    16'd18649: out <= 16'h07A3;    16'd18650: out <= 16'h04E2;    16'd18651: out <= 16'hFBFA;
    16'd18652: out <= 16'hFCE4;    16'd18653: out <= 16'h017C;    16'd18654: out <= 16'h0059;    16'd18655: out <= 16'h008A;
    16'd18656: out <= 16'h0206;    16'd18657: out <= 16'h0165;    16'd18658: out <= 16'h02DE;    16'd18659: out <= 16'hFEE5;
    16'd18660: out <= 16'hFF89;    16'd18661: out <= 16'hFF3C;    16'd18662: out <= 16'hFC34;    16'd18663: out <= 16'hF8B8;
    16'd18664: out <= 16'hFFA8;    16'd18665: out <= 16'h006F;    16'd18666: out <= 16'hFF69;    16'd18667: out <= 16'hFF2E;
    16'd18668: out <= 16'h0781;    16'd18669: out <= 16'hFDC1;    16'd18670: out <= 16'h03A4;    16'd18671: out <= 16'h02F3;
    16'd18672: out <= 16'hFE21;    16'd18673: out <= 16'hFDBD;    16'd18674: out <= 16'hFA6C;    16'd18675: out <= 16'h09E4;
    16'd18676: out <= 16'h0091;    16'd18677: out <= 16'hFFF9;    16'd18678: out <= 16'hFCB4;    16'd18679: out <= 16'hF57A;
    16'd18680: out <= 16'hFF5F;    16'd18681: out <= 16'hFE15;    16'd18682: out <= 16'hFA89;    16'd18683: out <= 16'h0304;
    16'd18684: out <= 16'h00CD;    16'd18685: out <= 16'hFE1D;    16'd18686: out <= 16'hFB69;    16'd18687: out <= 16'h0035;
    16'd18688: out <= 16'hFD96;    16'd18689: out <= 16'h06B4;    16'd18690: out <= 16'hFAEE;    16'd18691: out <= 16'h05C2;
    16'd18692: out <= 16'hFC43;    16'd18693: out <= 16'h024C;    16'd18694: out <= 16'h011F;    16'd18695: out <= 16'hFFEE;
    16'd18696: out <= 16'hFDAA;    16'd18697: out <= 16'hFFF5;    16'd18698: out <= 16'hFDA0;    16'd18699: out <= 16'hFEB3;
    16'd18700: out <= 16'hFE53;    16'd18701: out <= 16'h0120;    16'd18702: out <= 16'h0236;    16'd18703: out <= 16'h03F5;
    16'd18704: out <= 16'hF6F5;    16'd18705: out <= 16'h0402;    16'd18706: out <= 16'h0291;    16'd18707: out <= 16'h0280;
    16'd18708: out <= 16'h0876;    16'd18709: out <= 16'h0441;    16'd18710: out <= 16'h00BF;    16'd18711: out <= 16'hFD77;
    16'd18712: out <= 16'h0A52;    16'd18713: out <= 16'hFEA2;    16'd18714: out <= 16'hF9E8;    16'd18715: out <= 16'h0714;
    16'd18716: out <= 16'h0516;    16'd18717: out <= 16'h0686;    16'd18718: out <= 16'h080A;    16'd18719: out <= 16'h05CF;
    16'd18720: out <= 16'h00DD;    16'd18721: out <= 16'h03DB;    16'd18722: out <= 16'h0639;    16'd18723: out <= 16'h003E;
    16'd18724: out <= 16'h01A8;    16'd18725: out <= 16'hFF28;    16'd18726: out <= 16'h0843;    16'd18727: out <= 16'hFF95;
    16'd18728: out <= 16'h0714;    16'd18729: out <= 16'h0589;    16'd18730: out <= 16'h00D7;    16'd18731: out <= 16'h0324;
    16'd18732: out <= 16'hFE70;    16'd18733: out <= 16'h086C;    16'd18734: out <= 16'h0484;    16'd18735: out <= 16'hFCB4;
    16'd18736: out <= 16'h0050;    16'd18737: out <= 16'h03FC;    16'd18738: out <= 16'h0537;    16'd18739: out <= 16'h00EF;
    16'd18740: out <= 16'h03DB;    16'd18741: out <= 16'h04A1;    16'd18742: out <= 16'h0CA7;    16'd18743: out <= 16'h0AC3;
    16'd18744: out <= 16'h0682;    16'd18745: out <= 16'h0970;    16'd18746: out <= 16'h00D1;    16'd18747: out <= 16'h04A4;
    16'd18748: out <= 16'h0795;    16'd18749: out <= 16'h0726;    16'd18750: out <= 16'hFD34;    16'd18751: out <= 16'h03CD;
    16'd18752: out <= 16'h0845;    16'd18753: out <= 16'h00A7;    16'd18754: out <= 16'h020B;    16'd18755: out <= 16'h05EF;
    16'd18756: out <= 16'h0A13;    16'd18757: out <= 16'h0008;    16'd18758: out <= 16'h0175;    16'd18759: out <= 16'h00D2;
    16'd18760: out <= 16'h05EB;    16'd18761: out <= 16'h05C3;    16'd18762: out <= 16'h06DF;    16'd18763: out <= 16'hFD49;
    16'd18764: out <= 16'h04CD;    16'd18765: out <= 16'h027C;    16'd18766: out <= 16'h0223;    16'd18767: out <= 16'hFFE2;
    16'd18768: out <= 16'h01A4;    16'd18769: out <= 16'h0400;    16'd18770: out <= 16'h0051;    16'd18771: out <= 16'h03AE;
    16'd18772: out <= 16'h04CF;    16'd18773: out <= 16'h0679;    16'd18774: out <= 16'h042C;    16'd18775: out <= 16'h05AC;
    16'd18776: out <= 16'hFF5A;    16'd18777: out <= 16'h068F;    16'd18778: out <= 16'h0AAC;    16'd18779: out <= 16'h02E5;
    16'd18780: out <= 16'h0528;    16'd18781: out <= 16'h031E;    16'd18782: out <= 16'h03B3;    16'd18783: out <= 16'h04B4;
    16'd18784: out <= 16'h05C8;    16'd18785: out <= 16'h02AC;    16'd18786: out <= 16'h020B;    16'd18787: out <= 16'h0007;
    16'd18788: out <= 16'h049C;    16'd18789: out <= 16'h031D;    16'd18790: out <= 16'h023D;    16'd18791: out <= 16'h038D;
    16'd18792: out <= 16'h0AEC;    16'd18793: out <= 16'hFDAB;    16'd18794: out <= 16'h01C7;    16'd18795: out <= 16'hFA53;
    16'd18796: out <= 16'h06D5;    16'd18797: out <= 16'hFE1C;    16'd18798: out <= 16'h04E4;    16'd18799: out <= 16'h0805;
    16'd18800: out <= 16'h0342;    16'd18801: out <= 16'h0206;    16'd18802: out <= 16'h00BE;    16'd18803: out <= 16'hFEA5;
    16'd18804: out <= 16'h063C;    16'd18805: out <= 16'h0624;    16'd18806: out <= 16'hFEC9;    16'd18807: out <= 16'hFC49;
    16'd18808: out <= 16'h0133;    16'd18809: out <= 16'hFE93;    16'd18810: out <= 16'h08F3;    16'd18811: out <= 16'h0248;
    16'd18812: out <= 16'h00B1;    16'd18813: out <= 16'h0605;    16'd18814: out <= 16'h0466;    16'd18815: out <= 16'h070D;
    16'd18816: out <= 16'h0112;    16'd18817: out <= 16'h04DD;    16'd18818: out <= 16'h007C;    16'd18819: out <= 16'h04FE;
    16'd18820: out <= 16'h0717;    16'd18821: out <= 16'h0372;    16'd18822: out <= 16'hFD16;    16'd18823: out <= 16'h04BD;
    16'd18824: out <= 16'h013D;    16'd18825: out <= 16'h0636;    16'd18826: out <= 16'h02A3;    16'd18827: out <= 16'h0660;
    16'd18828: out <= 16'h040A;    16'd18829: out <= 16'h0402;    16'd18830: out <= 16'h0129;    16'd18831: out <= 16'h0798;
    16'd18832: out <= 16'h07E9;    16'd18833: out <= 16'h05AB;    16'd18834: out <= 16'h06F0;    16'd18835: out <= 16'h00C4;
    16'd18836: out <= 16'h01E2;    16'd18837: out <= 16'h046B;    16'd18838: out <= 16'hF696;    16'd18839: out <= 16'h06A0;
    16'd18840: out <= 16'h0761;    16'd18841: out <= 16'h0274;    16'd18842: out <= 16'h0307;    16'd18843: out <= 16'h0ACD;
    16'd18844: out <= 16'h019B;    16'd18845: out <= 16'h0804;    16'd18846: out <= 16'h0AA6;    16'd18847: out <= 16'h082E;
    16'd18848: out <= 16'h0664;    16'd18849: out <= 16'h052E;    16'd18850: out <= 16'h07A6;    16'd18851: out <= 16'h023F;
    16'd18852: out <= 16'hFC50;    16'd18853: out <= 16'h0B19;    16'd18854: out <= 16'h03E7;    16'd18855: out <= 16'h01C3;
    16'd18856: out <= 16'hFEE5;    16'd18857: out <= 16'h0137;    16'd18858: out <= 16'h0103;    16'd18859: out <= 16'h0465;
    16'd18860: out <= 16'h0881;    16'd18861: out <= 16'hFB77;    16'd18862: out <= 16'h0057;    16'd18863: out <= 16'h05C4;
    16'd18864: out <= 16'h0A77;    16'd18865: out <= 16'h0145;    16'd18866: out <= 16'h04E9;    16'd18867: out <= 16'h0578;
    16'd18868: out <= 16'h06C6;    16'd18869: out <= 16'h00B8;    16'd18870: out <= 16'h050B;    16'd18871: out <= 16'h0438;
    16'd18872: out <= 16'h0857;    16'd18873: out <= 16'h0612;    16'd18874: out <= 16'hFADA;    16'd18875: out <= 16'hFE61;
    16'd18876: out <= 16'h04A3;    16'd18877: out <= 16'hFFF9;    16'd18878: out <= 16'hFF58;    16'd18879: out <= 16'h0627;
    16'd18880: out <= 16'h009B;    16'd18881: out <= 16'h05EA;    16'd18882: out <= 16'h0162;    16'd18883: out <= 16'hFCB5;
    16'd18884: out <= 16'h01F0;    16'd18885: out <= 16'h0335;    16'd18886: out <= 16'h089A;    16'd18887: out <= 16'hFF06;
    16'd18888: out <= 16'h0C00;    16'd18889: out <= 16'h05AE;    16'd18890: out <= 16'h037B;    16'd18891: out <= 16'h07E6;
    16'd18892: out <= 16'h0578;    16'd18893: out <= 16'h0576;    16'd18894: out <= 16'h0262;    16'd18895: out <= 16'h0771;
    16'd18896: out <= 16'h01CD;    16'd18897: out <= 16'h008C;    16'd18898: out <= 16'h0A77;    16'd18899: out <= 16'h07F7;
    16'd18900: out <= 16'h00C3;    16'd18901: out <= 16'h0473;    16'd18902: out <= 16'h0476;    16'd18903: out <= 16'h08AA;
    16'd18904: out <= 16'hFD49;    16'd18905: out <= 16'h0367;    16'd18906: out <= 16'hF94F;    16'd18907: out <= 16'h001F;
    16'd18908: out <= 16'hFE1A;    16'd18909: out <= 16'h07DB;    16'd18910: out <= 16'hFDEF;    16'd18911: out <= 16'h04AA;
    16'd18912: out <= 16'hFC33;    16'd18913: out <= 16'hFFD8;    16'd18914: out <= 16'hFD30;    16'd18915: out <= 16'h02C5;
    16'd18916: out <= 16'hFA2E;    16'd18917: out <= 16'h003B;    16'd18918: out <= 16'hFD84;    16'd18919: out <= 16'h0203;
    16'd18920: out <= 16'hFF15;    16'd18921: out <= 16'h050A;    16'd18922: out <= 16'hFC96;    16'd18923: out <= 16'h003E;
    16'd18924: out <= 16'hFF4C;    16'd18925: out <= 16'hFE57;    16'd18926: out <= 16'hFF5C;    16'd18927: out <= 16'h0558;
    16'd18928: out <= 16'h0510;    16'd18929: out <= 16'h0009;    16'd18930: out <= 16'h0388;    16'd18931: out <= 16'hFBD3;
    16'd18932: out <= 16'h03CB;    16'd18933: out <= 16'hFB8A;    16'd18934: out <= 16'hFEE7;    16'd18935: out <= 16'h012C;
    16'd18936: out <= 16'h01F0;    16'd18937: out <= 16'hFDA8;    16'd18938: out <= 16'hFB83;    16'd18939: out <= 16'h0071;
    16'd18940: out <= 16'h0310;    16'd18941: out <= 16'hF7EA;    16'd18942: out <= 16'hFE73;    16'd18943: out <= 16'hFD44;
    16'd18944: out <= 16'h028C;    16'd18945: out <= 16'h0168;    16'd18946: out <= 16'hFDFE;    16'd18947: out <= 16'h04D2;
    16'd18948: out <= 16'hFE9B;    16'd18949: out <= 16'hFD37;    16'd18950: out <= 16'hF6F3;    16'd18951: out <= 16'hFDFB;
    16'd18952: out <= 16'hFDB1;    16'd18953: out <= 16'hFE01;    16'd18954: out <= 16'hFE95;    16'd18955: out <= 16'h0092;
    16'd18956: out <= 16'hFA40;    16'd18957: out <= 16'hFF0D;    16'd18958: out <= 16'h005E;    16'd18959: out <= 16'hFDFA;
    16'd18960: out <= 16'hFF1B;    16'd18961: out <= 16'h0165;    16'd18962: out <= 16'h00C9;    16'd18963: out <= 16'h0100;
    16'd18964: out <= 16'h03BF;    16'd18965: out <= 16'hFF5E;    16'd18966: out <= 16'hFFEF;    16'd18967: out <= 16'hFFCB;
    16'd18968: out <= 16'hFAA5;    16'd18969: out <= 16'hFFB1;    16'd18970: out <= 16'h011B;    16'd18971: out <= 16'h0428;
    16'd18972: out <= 16'h05CA;    16'd18973: out <= 16'h0387;    16'd18974: out <= 16'h034D;    16'd18975: out <= 16'h01EA;
    16'd18976: out <= 16'h0491;    16'd18977: out <= 16'h0598;    16'd18978: out <= 16'h0369;    16'd18979: out <= 16'h034E;
    16'd18980: out <= 16'h0711;    16'd18981: out <= 16'hFCF7;    16'd18982: out <= 16'h0BEA;    16'd18983: out <= 16'h0B06;
    16'd18984: out <= 16'h014E;    16'd18985: out <= 16'h03CF;    16'd18986: out <= 16'hF82C;    16'd18987: out <= 16'h06E9;
    16'd18988: out <= 16'h0B20;    16'd18989: out <= 16'h02A9;    16'd18990: out <= 16'h03D9;    16'd18991: out <= 16'h048C;
    16'd18992: out <= 16'hFFF0;    16'd18993: out <= 16'h08AD;    16'd18994: out <= 16'h010E;    16'd18995: out <= 16'h0064;
    16'd18996: out <= 16'h0267;    16'd18997: out <= 16'h061C;    16'd18998: out <= 16'hFBD3;    16'd18999: out <= 16'h024B;
    16'd19000: out <= 16'h00CF;    16'd19001: out <= 16'h05F9;    16'd19002: out <= 16'h0503;    16'd19003: out <= 16'hFE86;
    16'd19004: out <= 16'hFFED;    16'd19005: out <= 16'h07F0;    16'd19006: out <= 16'h052A;    16'd19007: out <= 16'h0D0B;
    16'd19008: out <= 16'h0ACA;    16'd19009: out <= 16'h0C7B;    16'd19010: out <= 16'hFE8C;    16'd19011: out <= 16'h00FE;
    16'd19012: out <= 16'h04E4;    16'd19013: out <= 16'h04CE;    16'd19014: out <= 16'hFF5D;    16'd19015: out <= 16'h0420;
    16'd19016: out <= 16'h0006;    16'd19017: out <= 16'h049D;    16'd19018: out <= 16'hFE08;    16'd19019: out <= 16'hFF94;
    16'd19020: out <= 16'h0212;    16'd19021: out <= 16'hFE9A;    16'd19022: out <= 16'h0388;    16'd19023: out <= 16'h0516;
    16'd19024: out <= 16'h06D2;    16'd19025: out <= 16'h060E;    16'd19026: out <= 16'hFFE4;    16'd19027: out <= 16'h0936;
    16'd19028: out <= 16'hFF5A;    16'd19029: out <= 16'h05DC;    16'd19030: out <= 16'h076A;    16'd19031: out <= 16'h0369;
    16'd19032: out <= 16'h03A5;    16'd19033: out <= 16'h0159;    16'd19034: out <= 16'h0B37;    16'd19035: out <= 16'h0185;
    16'd19036: out <= 16'h093B;    16'd19037: out <= 16'h044A;    16'd19038: out <= 16'h0143;    16'd19039: out <= 16'h02AB;
    16'd19040: out <= 16'h0500;    16'd19041: out <= 16'h075F;    16'd19042: out <= 16'h055F;    16'd19043: out <= 16'h0692;
    16'd19044: out <= 16'hFFA7;    16'd19045: out <= 16'hFF8C;    16'd19046: out <= 16'hFAE9;    16'd19047: out <= 16'h009D;
    16'd19048: out <= 16'h00B0;    16'd19049: out <= 16'h0151;    16'd19050: out <= 16'h005E;    16'd19051: out <= 16'hFE7D;
    16'd19052: out <= 16'h035F;    16'd19053: out <= 16'h07A2;    16'd19054: out <= 16'h0675;    16'd19055: out <= 16'h00FD;
    16'd19056: out <= 16'h0815;    16'd19057: out <= 16'h07A5;    16'd19058: out <= 16'hFFFD;    16'd19059: out <= 16'h032C;
    16'd19060: out <= 16'h0A5E;    16'd19061: out <= 16'h0715;    16'd19062: out <= 16'h01C4;    16'd19063: out <= 16'h0B9B;
    16'd19064: out <= 16'h0138;    16'd19065: out <= 16'h0078;    16'd19066: out <= 16'hFEAE;    16'd19067: out <= 16'h072E;
    16'd19068: out <= 16'h03FD;    16'd19069: out <= 16'hFFC6;    16'd19070: out <= 16'h0416;    16'd19071: out <= 16'h0343;
    16'd19072: out <= 16'h067C;    16'd19073: out <= 16'h0186;    16'd19074: out <= 16'h054B;    16'd19075: out <= 16'h0733;
    16'd19076: out <= 16'hFB18;    16'd19077: out <= 16'hFD7B;    16'd19078: out <= 16'h01CD;    16'd19079: out <= 16'h0082;
    16'd19080: out <= 16'h0314;    16'd19081: out <= 16'h00E1;    16'd19082: out <= 16'h0671;    16'd19083: out <= 16'h0A91;
    16'd19084: out <= 16'h0CD4;    16'd19085: out <= 16'h03A1;    16'd19086: out <= 16'h0484;    16'd19087: out <= 16'h03D5;
    16'd19088: out <= 16'h0C56;    16'd19089: out <= 16'hFE11;    16'd19090: out <= 16'hFF82;    16'd19091: out <= 16'h00D4;
    16'd19092: out <= 16'hFCD2;    16'd19093: out <= 16'h032C;    16'd19094: out <= 16'h03A5;    16'd19095: out <= 16'h0441;
    16'd19096: out <= 16'h0A91;    16'd19097: out <= 16'hFFB7;    16'd19098: out <= 16'h0201;    16'd19099: out <= 16'h0B96;
    16'd19100: out <= 16'h02F2;    16'd19101: out <= 16'h09B6;    16'd19102: out <= 16'h0BD2;    16'd19103: out <= 16'h0329;
    16'd19104: out <= 16'h138C;    16'd19105: out <= 16'h08D0;    16'd19106: out <= 16'h0311;    16'd19107: out <= 16'h049B;
    16'd19108: out <= 16'h00F9;    16'd19109: out <= 16'h0810;    16'd19110: out <= 16'h0159;    16'd19111: out <= 16'h0877;
    16'd19112: out <= 16'h03DB;    16'd19113: out <= 16'h02BF;    16'd19114: out <= 16'hFD73;    16'd19115: out <= 16'h01BD;
    16'd19116: out <= 16'h0626;    16'd19117: out <= 16'h06FC;    16'd19118: out <= 16'hFFF0;    16'd19119: out <= 16'h08D3;
    16'd19120: out <= 16'hFEBE;    16'd19121: out <= 16'hFBD6;    16'd19122: out <= 16'h00B9;    16'd19123: out <= 16'h03AC;
    16'd19124: out <= 16'hFFBC;    16'd19125: out <= 16'hFFF5;    16'd19126: out <= 16'h02D9;    16'd19127: out <= 16'h0659;
    16'd19128: out <= 16'h00D7;    16'd19129: out <= 16'h06A8;    16'd19130: out <= 16'h056F;    16'd19131: out <= 16'h04FD;
    16'd19132: out <= 16'h07B0;    16'd19133: out <= 16'hFE4E;    16'd19134: out <= 16'h05BC;    16'd19135: out <= 16'h03E4;
    16'd19136: out <= 16'h07C9;    16'd19137: out <= 16'h0273;    16'd19138: out <= 16'h02D0;    16'd19139: out <= 16'h0761;
    16'd19140: out <= 16'h0273;    16'd19141: out <= 16'h029B;    16'd19142: out <= 16'h01F6;    16'd19143: out <= 16'hFF29;
    16'd19144: out <= 16'h02D6;    16'd19145: out <= 16'h006D;    16'd19146: out <= 16'h03BA;    16'd19147: out <= 16'h068E;
    16'd19148: out <= 16'h01CD;    16'd19149: out <= 16'h01AB;    16'd19150: out <= 16'h028E;    16'd19151: out <= 16'h01FD;
    16'd19152: out <= 16'h008A;    16'd19153: out <= 16'h0808;    16'd19154: out <= 16'h0641;    16'd19155: out <= 16'h060A;
    16'd19156: out <= 16'h06FE;    16'd19157: out <= 16'h0715;    16'd19158: out <= 16'hFFA5;    16'd19159: out <= 16'h0536;
    16'd19160: out <= 16'h0934;    16'd19161: out <= 16'h0A50;    16'd19162: out <= 16'hFE83;    16'd19163: out <= 16'h0698;
    16'd19164: out <= 16'h0243;    16'd19165: out <= 16'h02C2;    16'd19166: out <= 16'h056B;    16'd19167: out <= 16'hFB22;
    16'd19168: out <= 16'hFC91;    16'd19169: out <= 16'hFFBF;    16'd19170: out <= 16'h0425;    16'd19171: out <= 16'hF994;
    16'd19172: out <= 16'hFCB0;    16'd19173: out <= 16'h0122;    16'd19174: out <= 16'hF933;    16'd19175: out <= 16'h07D9;
    16'd19176: out <= 16'hFDA5;    16'd19177: out <= 16'h0547;    16'd19178: out <= 16'hFBE2;    16'd19179: out <= 16'hFE8D;
    16'd19180: out <= 16'h0132;    16'd19181: out <= 16'hFF05;    16'd19182: out <= 16'h03E4;    16'd19183: out <= 16'hFFB8;
    16'd19184: out <= 16'hFDF9;    16'd19185: out <= 16'h0331;    16'd19186: out <= 16'h0364;    16'd19187: out <= 16'hFDB4;
    16'd19188: out <= 16'h01D8;    16'd19189: out <= 16'h00BB;    16'd19190: out <= 16'hFF16;    16'd19191: out <= 16'hF8A0;
    16'd19192: out <= 16'h0782;    16'd19193: out <= 16'h0553;    16'd19194: out <= 16'hF95E;    16'd19195: out <= 16'h03CE;
    16'd19196: out <= 16'hFB9F;    16'd19197: out <= 16'hF909;    16'd19198: out <= 16'hFF95;    16'd19199: out <= 16'hFF4C;
    16'd19200: out <= 16'h018E;    16'd19201: out <= 16'h07EB;    16'd19202: out <= 16'hFE56;    16'd19203: out <= 16'h0215;
    16'd19204: out <= 16'h0244;    16'd19205: out <= 16'hFE45;    16'd19206: out <= 16'hF747;    16'd19207: out <= 16'hFB85;
    16'd19208: out <= 16'hFB49;    16'd19209: out <= 16'h0534;    16'd19210: out <= 16'hFBAE;    16'd19211: out <= 16'hFFD2;
    16'd19212: out <= 16'h0034;    16'd19213: out <= 16'hFB57;    16'd19214: out <= 16'hFD55;    16'd19215: out <= 16'h00A5;
    16'd19216: out <= 16'h00ED;    16'd19217: out <= 16'hFDA9;    16'd19218: out <= 16'h0030;    16'd19219: out <= 16'h01AD;
    16'd19220: out <= 16'hFEA2;    16'd19221: out <= 16'h0345;    16'd19222: out <= 16'hF8B3;    16'd19223: out <= 16'h0745;
    16'd19224: out <= 16'hFAA2;    16'd19225: out <= 16'h0212;    16'd19226: out <= 16'h0152;    16'd19227: out <= 16'h045C;
    16'd19228: out <= 16'h0464;    16'd19229: out <= 16'hFD00;    16'd19230: out <= 16'h0347;    16'd19231: out <= 16'h018E;
    16'd19232: out <= 16'hFCB9;    16'd19233: out <= 16'h010A;    16'd19234: out <= 16'h0389;    16'd19235: out <= 16'h0293;
    16'd19236: out <= 16'h0030;    16'd19237: out <= 16'h05D6;    16'd19238: out <= 16'h05AB;    16'd19239: out <= 16'h03B6;
    16'd19240: out <= 16'h072C;    16'd19241: out <= 16'h02B4;    16'd19242: out <= 16'h07E6;    16'd19243: out <= 16'h02C5;
    16'd19244: out <= 16'hFF19;    16'd19245: out <= 16'h030B;    16'd19246: out <= 16'h0788;    16'd19247: out <= 16'h056B;
    16'd19248: out <= 16'hFFCE;    16'd19249: out <= 16'h0800;    16'd19250: out <= 16'h0895;    16'd19251: out <= 16'hFF88;
    16'd19252: out <= 16'h0010;    16'd19253: out <= 16'hFCBA;    16'd19254: out <= 16'h09C7;    16'd19255: out <= 16'hFE64;
    16'd19256: out <= 16'h0571;    16'd19257: out <= 16'h0618;    16'd19258: out <= 16'h0B45;    16'd19259: out <= 16'h0BB7;
    16'd19260: out <= 16'hF761;    16'd19261: out <= 16'h0597;    16'd19262: out <= 16'h00DA;    16'd19263: out <= 16'h0868;
    16'd19264: out <= 16'h0670;    16'd19265: out <= 16'hFFD8;    16'd19266: out <= 16'hFEDD;    16'd19267: out <= 16'hFF10;
    16'd19268: out <= 16'hFFA5;    16'd19269: out <= 16'h00FB;    16'd19270: out <= 16'h0349;    16'd19271: out <= 16'h09C1;
    16'd19272: out <= 16'hFC74;    16'd19273: out <= 16'h031A;    16'd19274: out <= 16'h024B;    16'd19275: out <= 16'h00B6;
    16'd19276: out <= 16'hFEF1;    16'd19277: out <= 16'h03E0;    16'd19278: out <= 16'h0241;    16'd19279: out <= 16'hFFDC;
    16'd19280: out <= 16'h0370;    16'd19281: out <= 16'h0579;    16'd19282: out <= 16'h0479;    16'd19283: out <= 16'h056D;
    16'd19284: out <= 16'h0173;    16'd19285: out <= 16'h0706;    16'd19286: out <= 16'h03E2;    16'd19287: out <= 16'hFF73;
    16'd19288: out <= 16'hFB9C;    16'd19289: out <= 16'h0385;    16'd19290: out <= 16'h09A3;    16'd19291: out <= 16'h0715;
    16'd19292: out <= 16'h048D;    16'd19293: out <= 16'h0243;    16'd19294: out <= 16'hFF7B;    16'd19295: out <= 16'h07E5;
    16'd19296: out <= 16'h005C;    16'd19297: out <= 16'h060C;    16'd19298: out <= 16'h02D8;    16'd19299: out <= 16'h02EE;
    16'd19300: out <= 16'h07E0;    16'd19301: out <= 16'h0211;    16'd19302: out <= 16'h0855;    16'd19303: out <= 16'h0713;
    16'd19304: out <= 16'h0059;    16'd19305: out <= 16'h05CC;    16'd19306: out <= 16'h071E;    16'd19307: out <= 16'h033A;
    16'd19308: out <= 16'h026B;    16'd19309: out <= 16'h02E2;    16'd19310: out <= 16'h006F;    16'd19311: out <= 16'hFD30;
    16'd19312: out <= 16'hFEC6;    16'd19313: out <= 16'h03D3;    16'd19314: out <= 16'h00C6;    16'd19315: out <= 16'h01B9;
    16'd19316: out <= 16'h00A6;    16'd19317: out <= 16'h02D8;    16'd19318: out <= 16'hFC52;    16'd19319: out <= 16'h0601;
    16'd19320: out <= 16'h0334;    16'd19321: out <= 16'h009E;    16'd19322: out <= 16'h0824;    16'd19323: out <= 16'hFF35;
    16'd19324: out <= 16'h0622;    16'd19325: out <= 16'h08F5;    16'd19326: out <= 16'h0462;    16'd19327: out <= 16'hFC3C;
    16'd19328: out <= 16'h0441;    16'd19329: out <= 16'h0A15;    16'd19330: out <= 16'h0465;    16'd19331: out <= 16'hFFDA;
    16'd19332: out <= 16'hFD46;    16'd19333: out <= 16'h0089;    16'd19334: out <= 16'h038C;    16'd19335: out <= 16'h035B;
    16'd19336: out <= 16'h0243;    16'd19337: out <= 16'h0401;    16'd19338: out <= 16'h068C;    16'd19339: out <= 16'hFA71;
    16'd19340: out <= 16'h09E7;    16'd19341: out <= 16'h0A0A;    16'd19342: out <= 16'h02FD;    16'd19343: out <= 16'h0475;
    16'd19344: out <= 16'h01D1;    16'd19345: out <= 16'h0658;    16'd19346: out <= 16'h0A73;    16'd19347: out <= 16'h0537;
    16'd19348: out <= 16'h03AF;    16'd19349: out <= 16'hFABD;    16'd19350: out <= 16'h07BF;    16'd19351: out <= 16'hFD50;
    16'd19352: out <= 16'h050B;    16'd19353: out <= 16'h05A8;    16'd19354: out <= 16'hFFCF;    16'd19355: out <= 16'hFF54;
    16'd19356: out <= 16'h0299;    16'd19357: out <= 16'hFF83;    16'd19358: out <= 16'h0565;    16'd19359: out <= 16'h018E;
    16'd19360: out <= 16'h046F;    16'd19361: out <= 16'h01F9;    16'd19362: out <= 16'h06C0;    16'd19363: out <= 16'h03B6;
    16'd19364: out <= 16'h0543;    16'd19365: out <= 16'h02CB;    16'd19366: out <= 16'hFC44;    16'd19367: out <= 16'h0923;
    16'd19368: out <= 16'h027A;    16'd19369: out <= 16'h004F;    16'd19370: out <= 16'h00F1;    16'd19371: out <= 16'h01BE;
    16'd19372: out <= 16'h0352;    16'd19373: out <= 16'h0635;    16'd19374: out <= 16'h0979;    16'd19375: out <= 16'h0BF2;
    16'd19376: out <= 16'h05AF;    16'd19377: out <= 16'h050A;    16'd19378: out <= 16'h00E7;    16'd19379: out <= 16'h04B0;
    16'd19380: out <= 16'h03A1;    16'd19381: out <= 16'h00CD;    16'd19382: out <= 16'hF9A2;    16'd19383: out <= 16'h03D1;
    16'd19384: out <= 16'h073B;    16'd19385: out <= 16'h0527;    16'd19386: out <= 16'h0010;    16'd19387: out <= 16'h058F;
    16'd19388: out <= 16'h02F7;    16'd19389: out <= 16'h07E2;    16'd19390: out <= 16'h0444;    16'd19391: out <= 16'h0897;
    16'd19392: out <= 16'h00D3;    16'd19393: out <= 16'h0727;    16'd19394: out <= 16'hFC75;    16'd19395: out <= 16'h04F7;
    16'd19396: out <= 16'h02E8;    16'd19397: out <= 16'h0A53;    16'd19398: out <= 16'h08CF;    16'd19399: out <= 16'h0ABA;
    16'd19400: out <= 16'h01B9;    16'd19401: out <= 16'h0111;    16'd19402: out <= 16'h040C;    16'd19403: out <= 16'h07A4;
    16'd19404: out <= 16'h0544;    16'd19405: out <= 16'h0007;    16'd19406: out <= 16'h0B1D;    16'd19407: out <= 16'h035A;
    16'd19408: out <= 16'hFF96;    16'd19409: out <= 16'h05C1;    16'd19410: out <= 16'hFEF5;    16'd19411: out <= 16'h0561;
    16'd19412: out <= 16'hFED3;    16'd19413: out <= 16'h0716;    16'd19414: out <= 16'h03C4;    16'd19415: out <= 16'h0348;
    16'd19416: out <= 16'h033B;    16'd19417: out <= 16'hF9A4;    16'd19418: out <= 16'h0067;    16'd19419: out <= 16'h0BDC;
    16'd19420: out <= 16'h01FD;    16'd19421: out <= 16'hFAA5;    16'd19422: out <= 16'hFD00;    16'd19423: out <= 16'h02B4;
    16'd19424: out <= 16'h0066;    16'd19425: out <= 16'h04DF;    16'd19426: out <= 16'h0603;    16'd19427: out <= 16'h004C;
    16'd19428: out <= 16'hFECD;    16'd19429: out <= 16'hFE5C;    16'd19430: out <= 16'h01DF;    16'd19431: out <= 16'h0154;
    16'd19432: out <= 16'h0505;    16'd19433: out <= 16'hFDCE;    16'd19434: out <= 16'h001E;    16'd19435: out <= 16'hFF4B;
    16'd19436: out <= 16'h0247;    16'd19437: out <= 16'hFFCE;    16'd19438: out <= 16'hFD7D;    16'd19439: out <= 16'hF89C;
    16'd19440: out <= 16'h00B1;    16'd19441: out <= 16'h01DB;    16'd19442: out <= 16'h017A;    16'd19443: out <= 16'h002E;
    16'd19444: out <= 16'hFE0D;    16'd19445: out <= 16'h0164;    16'd19446: out <= 16'h04BF;    16'd19447: out <= 16'hFD50;
    16'd19448: out <= 16'hFDF1;    16'd19449: out <= 16'hFEE9;    16'd19450: out <= 16'hFDF5;    16'd19451: out <= 16'hFF11;
    16'd19452: out <= 16'h002C;    16'd19453: out <= 16'h019B;    16'd19454: out <= 16'hFC36;    16'd19455: out <= 16'h0199;
    16'd19456: out <= 16'h080C;    16'd19457: out <= 16'hFE93;    16'd19458: out <= 16'hFF9D;    16'd19459: out <= 16'h018E;
    16'd19460: out <= 16'hFFDE;    16'd19461: out <= 16'h00A6;    16'd19462: out <= 16'hFF6B;    16'd19463: out <= 16'h038F;
    16'd19464: out <= 16'h0108;    16'd19465: out <= 16'hFB9F;    16'd19466: out <= 16'hFEB2;    16'd19467: out <= 16'hFE29;
    16'd19468: out <= 16'h0488;    16'd19469: out <= 16'hFD39;    16'd19470: out <= 16'h00DB;    16'd19471: out <= 16'hFCE0;
    16'd19472: out <= 16'h0463;    16'd19473: out <= 16'h0549;    16'd19474: out <= 16'hFBF1;    16'd19475: out <= 16'h049B;
    16'd19476: out <= 16'hFFEB;    16'd19477: out <= 16'h04FD;    16'd19478: out <= 16'hFDCC;    16'd19479: out <= 16'hFACC;
    16'd19480: out <= 16'h01AC;    16'd19481: out <= 16'h0153;    16'd19482: out <= 16'h05BB;    16'd19483: out <= 16'h0784;
    16'd19484: out <= 16'h03C9;    16'd19485: out <= 16'h05C9;    16'd19486: out <= 16'h0351;    16'd19487: out <= 16'h047A;
    16'd19488: out <= 16'h056D;    16'd19489: out <= 16'h0501;    16'd19490: out <= 16'h08C8;    16'd19491: out <= 16'h07A8;
    16'd19492: out <= 16'h0735;    16'd19493: out <= 16'hFFCD;    16'd19494: out <= 16'h0625;    16'd19495: out <= 16'h0AC1;
    16'd19496: out <= 16'h03A6;    16'd19497: out <= 16'hFDD1;    16'd19498: out <= 16'h09C7;    16'd19499: out <= 16'h03F2;
    16'd19500: out <= 16'h06CC;    16'd19501: out <= 16'h0800;    16'd19502: out <= 16'hFDFC;    16'd19503: out <= 16'h01D9;
    16'd19504: out <= 16'h00DB;    16'd19505: out <= 16'h0419;    16'd19506: out <= 16'h0066;    16'd19507: out <= 16'h003E;
    16'd19508: out <= 16'h0435;    16'd19509: out <= 16'h03E9;    16'd19510: out <= 16'h0153;    16'd19511: out <= 16'hFEDA;
    16'd19512: out <= 16'h059C;    16'd19513: out <= 16'h037B;    16'd19514: out <= 16'h005B;    16'd19515: out <= 16'h03DF;
    16'd19516: out <= 16'h040F;    16'd19517: out <= 16'h0ABB;    16'd19518: out <= 16'h011D;    16'd19519: out <= 16'h0720;
    16'd19520: out <= 16'h02EC;    16'd19521: out <= 16'h000E;    16'd19522: out <= 16'h000F;    16'd19523: out <= 16'hFA04;
    16'd19524: out <= 16'h07C0;    16'd19525: out <= 16'h05FD;    16'd19526: out <= 16'h0402;    16'd19527: out <= 16'h0375;
    16'd19528: out <= 16'h0431;    16'd19529: out <= 16'hFB1A;    16'd19530: out <= 16'h0CB0;    16'd19531: out <= 16'h02B2;
    16'd19532: out <= 16'h01F0;    16'd19533: out <= 16'h038B;    16'd19534: out <= 16'h0204;    16'd19535: out <= 16'h0646;
    16'd19536: out <= 16'h05F7;    16'd19537: out <= 16'h0433;    16'd19538: out <= 16'h04CB;    16'd19539: out <= 16'h034C;
    16'd19540: out <= 16'h01FC;    16'd19541: out <= 16'h048B;    16'd19542: out <= 16'h0308;    16'd19543: out <= 16'h0358;
    16'd19544: out <= 16'h0431;    16'd19545: out <= 16'h07AF;    16'd19546: out <= 16'h0854;    16'd19547: out <= 16'h0150;
    16'd19548: out <= 16'h031F;    16'd19549: out <= 16'h0209;    16'd19550: out <= 16'h0332;    16'd19551: out <= 16'h0622;
    16'd19552: out <= 16'h08A8;    16'd19553: out <= 16'h06BF;    16'd19554: out <= 16'h0982;    16'd19555: out <= 16'h05EF;
    16'd19556: out <= 16'hFC20;    16'd19557: out <= 16'h02F7;    16'd19558: out <= 16'h098C;    16'd19559: out <= 16'h02CD;
    16'd19560: out <= 16'hFD6A;    16'd19561: out <= 16'h0469;    16'd19562: out <= 16'hFD04;    16'd19563: out <= 16'h01F8;
    16'd19564: out <= 16'h0407;    16'd19565: out <= 16'hFF1D;    16'd19566: out <= 16'h0AAA;    16'd19567: out <= 16'h04D2;
    16'd19568: out <= 16'h09B7;    16'd19569: out <= 16'h0514;    16'd19570: out <= 16'hFD75;    16'd19571: out <= 16'h0231;
    16'd19572: out <= 16'h0274;    16'd19573: out <= 16'h05FE;    16'd19574: out <= 16'h049D;    16'd19575: out <= 16'h07E9;
    16'd19576: out <= 16'h05F8;    16'd19577: out <= 16'h073E;    16'd19578: out <= 16'h0301;    16'd19579: out <= 16'hF9E7;
    16'd19580: out <= 16'h071F;    16'd19581: out <= 16'hFF10;    16'd19582: out <= 16'hFF8E;    16'd19583: out <= 16'h039D;
    16'd19584: out <= 16'h085B;    16'd19585: out <= 16'h0346;    16'd19586: out <= 16'h027A;    16'd19587: out <= 16'h03F3;
    16'd19588: out <= 16'hFE90;    16'd19589: out <= 16'h0314;    16'd19590: out <= 16'h040B;    16'd19591: out <= 16'h0373;
    16'd19592: out <= 16'h0474;    16'd19593: out <= 16'h0168;    16'd19594: out <= 16'h0809;    16'd19595: out <= 16'h034A;
    16'd19596: out <= 16'h0A7A;    16'd19597: out <= 16'h03A1;    16'd19598: out <= 16'h05FE;    16'd19599: out <= 16'hFF76;
    16'd19600: out <= 16'h0CF6;    16'd19601: out <= 16'h0369;    16'd19602: out <= 16'h02D5;    16'd19603: out <= 16'h00FB;
    16'd19604: out <= 16'h0C7B;    16'd19605: out <= 16'h06A4;    16'd19606: out <= 16'h0185;    16'd19607: out <= 16'hFF28;
    16'd19608: out <= 16'h062F;    16'd19609: out <= 16'h044F;    16'd19610: out <= 16'h00A3;    16'd19611: out <= 16'hFCAD;
    16'd19612: out <= 16'h04B0;    16'd19613: out <= 16'h0847;    16'd19614: out <= 16'h081B;    16'd19615: out <= 16'h0217;
    16'd19616: out <= 16'h0971;    16'd19617: out <= 16'hFBDD;    16'd19618: out <= 16'h070A;    16'd19619: out <= 16'hFFEB;
    16'd19620: out <= 16'h0378;    16'd19621: out <= 16'hFF88;    16'd19622: out <= 16'h058B;    16'd19623: out <= 16'h0350;
    16'd19624: out <= 16'h00FF;    16'd19625: out <= 16'h0293;    16'd19626: out <= 16'h0533;    16'd19627: out <= 16'h032E;
    16'd19628: out <= 16'hFF2F;    16'd19629: out <= 16'hFAFC;    16'd19630: out <= 16'h070C;    16'd19631: out <= 16'h07F1;
    16'd19632: out <= 16'h0125;    16'd19633: out <= 16'h03A0;    16'd19634: out <= 16'h0029;    16'd19635: out <= 16'h0428;
    16'd19636: out <= 16'h0765;    16'd19637: out <= 16'h080E;    16'd19638: out <= 16'hFFF3;    16'd19639: out <= 16'h061B;
    16'd19640: out <= 16'h0502;    16'd19641: out <= 16'h0BD2;    16'd19642: out <= 16'hFF10;    16'd19643: out <= 16'h03A8;
    16'd19644: out <= 16'h0A06;    16'd19645: out <= 16'hFC65;    16'd19646: out <= 16'h051C;    16'd19647: out <= 16'h0402;
    16'd19648: out <= 16'hFFB4;    16'd19649: out <= 16'h0179;    16'd19650: out <= 16'h0A96;    16'd19651: out <= 16'hFCBA;
    16'd19652: out <= 16'h0309;    16'd19653: out <= 16'h056C;    16'd19654: out <= 16'h0194;    16'd19655: out <= 16'hFF82;
    16'd19656: out <= 16'h0005;    16'd19657: out <= 16'h036C;    16'd19658: out <= 16'h0279;    16'd19659: out <= 16'hFC93;
    16'd19660: out <= 16'hFB71;    16'd19661: out <= 16'hFD28;    16'd19662: out <= 16'hFEAE;    16'd19663: out <= 16'h01AE;
    16'd19664: out <= 16'h02E0;    16'd19665: out <= 16'h0605;    16'd19666: out <= 16'hFFB8;    16'd19667: out <= 16'h0440;
    16'd19668: out <= 16'hFF2E;    16'd19669: out <= 16'h05FC;    16'd19670: out <= 16'h055A;    16'd19671: out <= 16'h0738;
    16'd19672: out <= 16'hFB33;    16'd19673: out <= 16'hFC1E;    16'd19674: out <= 16'h04E7;    16'd19675: out <= 16'h0454;
    16'd19676: out <= 16'h094C;    16'd19677: out <= 16'hFA15;    16'd19678: out <= 16'hFFB4;    16'd19679: out <= 16'hFD0C;
    16'd19680: out <= 16'h03D0;    16'd19681: out <= 16'hFF93;    16'd19682: out <= 16'hFFE0;    16'd19683: out <= 16'h050D;
    16'd19684: out <= 16'h028F;    16'd19685: out <= 16'hFD25;    16'd19686: out <= 16'h0115;    16'd19687: out <= 16'hFB8A;
    16'd19688: out <= 16'h056E;    16'd19689: out <= 16'h055D;    16'd19690: out <= 16'hFD60;    16'd19691: out <= 16'h0053;
    16'd19692: out <= 16'h0082;    16'd19693: out <= 16'hFE2C;    16'd19694: out <= 16'h0B19;    16'd19695: out <= 16'h02AF;
    16'd19696: out <= 16'hFF3E;    16'd19697: out <= 16'hFD84;    16'd19698: out <= 16'hFAD4;    16'd19699: out <= 16'h01D3;
    16'd19700: out <= 16'hFF88;    16'd19701: out <= 16'hFFEE;    16'd19702: out <= 16'hFA71;    16'd19703: out <= 16'hFEA4;
    16'd19704: out <= 16'hFE26;    16'd19705: out <= 16'hFFE7;    16'd19706: out <= 16'hF9E6;    16'd19707: out <= 16'hFE43;
    16'd19708: out <= 16'h019F;    16'd19709: out <= 16'h0140;    16'd19710: out <= 16'hFF0C;    16'd19711: out <= 16'hFF29;
    16'd19712: out <= 16'h07A3;    16'd19713: out <= 16'h050F;    16'd19714: out <= 16'h0028;    16'd19715: out <= 16'h0584;
    16'd19716: out <= 16'h025F;    16'd19717: out <= 16'hFAEB;    16'd19718: out <= 16'hFCC8;    16'd19719: out <= 16'h009C;
    16'd19720: out <= 16'hFA78;    16'd19721: out <= 16'hFE82;    16'd19722: out <= 16'h0333;    16'd19723: out <= 16'h04C2;
    16'd19724: out <= 16'h0290;    16'd19725: out <= 16'hFF64;    16'd19726: out <= 16'h0178;    16'd19727: out <= 16'h0108;
    16'd19728: out <= 16'hF999;    16'd19729: out <= 16'h097A;    16'd19730: out <= 16'h00E8;    16'd19731: out <= 16'h05D6;
    16'd19732: out <= 16'hFFD6;    16'd19733: out <= 16'hFF1C;    16'd19734: out <= 16'h0027;    16'd19735: out <= 16'h00B7;
    16'd19736: out <= 16'hFAB2;    16'd19737: out <= 16'hFF06;    16'd19738: out <= 16'h00F2;    16'd19739: out <= 16'h077A;
    16'd19740: out <= 16'hFBED;    16'd19741: out <= 16'h04CD;    16'd19742: out <= 16'h025B;    16'd19743: out <= 16'h050F;
    16'd19744: out <= 16'h052A;    16'd19745: out <= 16'h03BE;    16'd19746: out <= 16'h0964;    16'd19747: out <= 16'h07DE;
    16'd19748: out <= 16'h053F;    16'd19749: out <= 16'h0AFA;    16'd19750: out <= 16'h0881;    16'd19751: out <= 16'hFE3D;
    16'd19752: out <= 16'h0305;    16'd19753: out <= 16'hFDE1;    16'd19754: out <= 16'h078D;    16'd19755: out <= 16'h06EF;
    16'd19756: out <= 16'hFDA8;    16'd19757: out <= 16'h0739;    16'd19758: out <= 16'hFC76;    16'd19759: out <= 16'h0089;
    16'd19760: out <= 16'h00EE;    16'd19761: out <= 16'h03F6;    16'd19762: out <= 16'h0A7E;    16'd19763: out <= 16'hFC94;
    16'd19764: out <= 16'h07EE;    16'd19765: out <= 16'h0586;    16'd19766: out <= 16'h08B3;    16'd19767: out <= 16'h00F6;
    16'd19768: out <= 16'h04DE;    16'd19769: out <= 16'h0789;    16'd19770: out <= 16'h02E4;    16'd19771: out <= 16'h0D60;
    16'd19772: out <= 16'h048D;    16'd19773: out <= 16'h022C;    16'd19774: out <= 16'h060C;    16'd19775: out <= 16'h01A1;
    16'd19776: out <= 16'h0314;    16'd19777: out <= 16'h090E;    16'd19778: out <= 16'h090C;    16'd19779: out <= 16'h01C0;
    16'd19780: out <= 16'h0324;    16'd19781: out <= 16'h03BD;    16'd19782: out <= 16'h0176;    16'd19783: out <= 16'hFFC4;
    16'd19784: out <= 16'h054F;    16'd19785: out <= 16'h0411;    16'd19786: out <= 16'h060B;    16'd19787: out <= 16'hFF61;
    16'd19788: out <= 16'h06B4;    16'd19789: out <= 16'hFECC;    16'd19790: out <= 16'h05DE;    16'd19791: out <= 16'h0173;
    16'd19792: out <= 16'h00CE;    16'd19793: out <= 16'h0405;    16'd19794: out <= 16'hFFC1;    16'd19795: out <= 16'h0186;
    16'd19796: out <= 16'h07C7;    16'd19797: out <= 16'h0136;    16'd19798: out <= 16'h056D;    16'd19799: out <= 16'h06F3;
    16'd19800: out <= 16'h0CAB;    16'd19801: out <= 16'h0A66;    16'd19802: out <= 16'h0515;    16'd19803: out <= 16'h017F;
    16'd19804: out <= 16'h08A1;    16'd19805: out <= 16'h07F4;    16'd19806: out <= 16'h099A;    16'd19807: out <= 16'h0B6E;
    16'd19808: out <= 16'h045C;    16'd19809: out <= 16'h051F;    16'd19810: out <= 16'h0450;    16'd19811: out <= 16'h0AAB;
    16'd19812: out <= 16'hFED0;    16'd19813: out <= 16'h05B4;    16'd19814: out <= 16'h07FA;    16'd19815: out <= 16'h0B77;
    16'd19816: out <= 16'h0549;    16'd19817: out <= 16'h020C;    16'd19818: out <= 16'h073D;    16'd19819: out <= 16'h00DD;
    16'd19820: out <= 16'h00F8;    16'd19821: out <= 16'h05FD;    16'd19822: out <= 16'h037A;    16'd19823: out <= 16'h033E;
    16'd19824: out <= 16'h0769;    16'd19825: out <= 16'h0410;    16'd19826: out <= 16'h0932;    16'd19827: out <= 16'hFFD6;
    16'd19828: out <= 16'h021C;    16'd19829: out <= 16'h0162;    16'd19830: out <= 16'h020A;    16'd19831: out <= 16'h0297;
    16'd19832: out <= 16'h082A;    16'd19833: out <= 16'hFD92;    16'd19834: out <= 16'h064C;    16'd19835: out <= 16'h0073;
    16'd19836: out <= 16'h04FF;    16'd19837: out <= 16'h0769;    16'd19838: out <= 16'h017F;    16'd19839: out <= 16'h039D;
    16'd19840: out <= 16'h000B;    16'd19841: out <= 16'h00B2;    16'd19842: out <= 16'h01BB;    16'd19843: out <= 16'h06C9;
    16'd19844: out <= 16'hFB97;    16'd19845: out <= 16'h04F2;    16'd19846: out <= 16'h0106;    16'd19847: out <= 16'h033D;
    16'd19848: out <= 16'hFF07;    16'd19849: out <= 16'h04C8;    16'd19850: out <= 16'h02B5;    16'd19851: out <= 16'h05A9;
    16'd19852: out <= 16'hFE23;    16'd19853: out <= 16'hFFA3;    16'd19854: out <= 16'hFF50;    16'd19855: out <= 16'h048A;
    16'd19856: out <= 16'hF8EF;    16'd19857: out <= 16'h01FE;    16'd19858: out <= 16'h0220;    16'd19859: out <= 16'h0374;
    16'd19860: out <= 16'h06F0;    16'd19861: out <= 16'hFDE2;    16'd19862: out <= 16'h0DB4;    16'd19863: out <= 16'hFDED;
    16'd19864: out <= 16'hFEC3;    16'd19865: out <= 16'h067B;    16'd19866: out <= 16'h05ED;    16'd19867: out <= 16'h029E;
    16'd19868: out <= 16'h05B9;    16'd19869: out <= 16'hFF6F;    16'd19870: out <= 16'h02BA;    16'd19871: out <= 16'hFD9D;
    16'd19872: out <= 16'hFDE7;    16'd19873: out <= 16'h041E;    16'd19874: out <= 16'h07F2;    16'd19875: out <= 16'hFEFE;
    16'd19876: out <= 16'h069A;    16'd19877: out <= 16'h030A;    16'd19878: out <= 16'h0264;    16'd19879: out <= 16'h00B3;
    16'd19880: out <= 16'h06C8;    16'd19881: out <= 16'h0473;    16'd19882: out <= 16'hFFA1;    16'd19883: out <= 16'h0021;
    16'd19884: out <= 16'h0390;    16'd19885: out <= 16'hFED4;    16'd19886: out <= 16'hFE1D;    16'd19887: out <= 16'h0716;
    16'd19888: out <= 16'h067E;    16'd19889: out <= 16'h0B3D;    16'd19890: out <= 16'h005C;    16'd19891: out <= 16'h062A;
    16'd19892: out <= 16'h040F;    16'd19893: out <= 16'h06C9;    16'd19894: out <= 16'h09BA;    16'd19895: out <= 16'h0363;
    16'd19896: out <= 16'h0114;    16'd19897: out <= 16'h0469;    16'd19898: out <= 16'h036F;    16'd19899: out <= 16'h0392;
    16'd19900: out <= 16'h023A;    16'd19901: out <= 16'hFF80;    16'd19902: out <= 16'h0A6E;    16'd19903: out <= 16'hFF6A;
    16'd19904: out <= 16'h04CE;    16'd19905: out <= 16'h0477;    16'd19906: out <= 16'h027C;    16'd19907: out <= 16'h0ACD;
    16'd19908: out <= 16'h026E;    16'd19909: out <= 16'hFE1B;    16'd19910: out <= 16'h00DF;    16'd19911: out <= 16'h0242;
    16'd19912: out <= 16'h0232;    16'd19913: out <= 16'h0818;    16'd19914: out <= 16'h0945;    16'd19915: out <= 16'h0483;
    16'd19916: out <= 16'h0415;    16'd19917: out <= 16'h04FB;    16'd19918: out <= 16'h02F2;    16'd19919: out <= 16'h02EF;
    16'd19920: out <= 16'h078A;    16'd19921: out <= 16'h0384;    16'd19922: out <= 16'h0011;    16'd19923: out <= 16'h092E;
    16'd19924: out <= 16'hF91B;    16'd19925: out <= 16'h04ED;    16'd19926: out <= 16'hFC65;    16'd19927: out <= 16'h07B5;
    16'd19928: out <= 16'h0AE5;    16'd19929: out <= 16'hFD85;    16'd19930: out <= 16'h03D1;    16'd19931: out <= 16'h06AE;
    16'd19932: out <= 16'hFD21;    16'd19933: out <= 16'hF914;    16'd19934: out <= 16'hFD33;    16'd19935: out <= 16'hFD90;
    16'd19936: out <= 16'hF798;    16'd19937: out <= 16'h0453;    16'd19938: out <= 16'h00E2;    16'd19939: out <= 16'hFA79;
    16'd19940: out <= 16'h0121;    16'd19941: out <= 16'h01B8;    16'd19942: out <= 16'h04B5;    16'd19943: out <= 16'h0564;
    16'd19944: out <= 16'h01EF;    16'd19945: out <= 16'h037B;    16'd19946: out <= 16'h0256;    16'd19947: out <= 16'hFA2C;
    16'd19948: out <= 16'hFB6B;    16'd19949: out <= 16'h0034;    16'd19950: out <= 16'hFD00;    16'd19951: out <= 16'hFD9C;
    16'd19952: out <= 16'h0411;    16'd19953: out <= 16'hFE1D;    16'd19954: out <= 16'hF9BE;    16'd19955: out <= 16'hFA01;
    16'd19956: out <= 16'h04DC;    16'd19957: out <= 16'hFF9E;    16'd19958: out <= 16'h046A;    16'd19959: out <= 16'h0371;
    16'd19960: out <= 16'hFDAC;    16'd19961: out <= 16'hF80C;    16'd19962: out <= 16'h03B3;    16'd19963: out <= 16'h02DB;
    16'd19964: out <= 16'h0239;    16'd19965: out <= 16'h01C8;    16'd19966: out <= 16'hF904;    16'd19967: out <= 16'hFCAF;
    16'd19968: out <= 16'h01D2;    16'd19969: out <= 16'hFEC5;    16'd19970: out <= 16'hFF45;    16'd19971: out <= 16'h023A;
    16'd19972: out <= 16'h026B;    16'd19973: out <= 16'h0160;    16'd19974: out <= 16'hFE54;    16'd19975: out <= 16'h0067;
    16'd19976: out <= 16'hFF6C;    16'd19977: out <= 16'hFABD;    16'd19978: out <= 16'h0485;    16'd19979: out <= 16'h0203;
    16'd19980: out <= 16'hFAAD;    16'd19981: out <= 16'h0185;    16'd19982: out <= 16'h0178;    16'd19983: out <= 16'h025B;
    16'd19984: out <= 16'h0451;    16'd19985: out <= 16'hFC9B;    16'd19986: out <= 16'h0258;    16'd19987: out <= 16'hFC82;
    16'd19988: out <= 16'hFC04;    16'd19989: out <= 16'h0332;    16'd19990: out <= 16'hFF87;    16'd19991: out <= 16'h0313;
    16'd19992: out <= 16'h0728;    16'd19993: out <= 16'hFA97;    16'd19994: out <= 16'h09D2;    16'd19995: out <= 16'h0DB2;
    16'd19996: out <= 16'h0417;    16'd19997: out <= 16'h03CF;    16'd19998: out <= 16'h055C;    16'd19999: out <= 16'h0205;
    16'd20000: out <= 16'hFDEE;    16'd20001: out <= 16'hF91E;    16'd20002: out <= 16'hFD7A;    16'd20003: out <= 16'hFF68;
    16'd20004: out <= 16'h051C;    16'd20005: out <= 16'h06D8;    16'd20006: out <= 16'h00E8;    16'd20007: out <= 16'h0AD9;
    16'd20008: out <= 16'h06BB;    16'd20009: out <= 16'h01E9;    16'd20010: out <= 16'h038D;    16'd20011: out <= 16'h01F9;
    16'd20012: out <= 16'h054B;    16'd20013: out <= 16'h0BD4;    16'd20014: out <= 16'h0494;    16'd20015: out <= 16'h00B3;
    16'd20016: out <= 16'h09D7;    16'd20017: out <= 16'h03E6;    16'd20018: out <= 16'h05D3;    16'd20019: out <= 16'h02C0;
    16'd20020: out <= 16'h0D57;    16'd20021: out <= 16'hFFE5;    16'd20022: out <= 16'h066E;    16'd20023: out <= 16'h0390;
    16'd20024: out <= 16'hFB98;    16'd20025: out <= 16'h036E;    16'd20026: out <= 16'h0633;    16'd20027: out <= 16'h07C3;
    16'd20028: out <= 16'h024E;    16'd20029: out <= 16'h0ADF;    16'd20030: out <= 16'h077F;    16'd20031: out <= 16'h028A;
    16'd20032: out <= 16'h0588;    16'd20033: out <= 16'h02B4;    16'd20034: out <= 16'h0A2A;    16'd20035: out <= 16'h0B34;
    16'd20036: out <= 16'h03EF;    16'd20037: out <= 16'h0412;    16'd20038: out <= 16'h04BE;    16'd20039: out <= 16'h0E3C;
    16'd20040: out <= 16'h06C7;    16'd20041: out <= 16'h070B;    16'd20042: out <= 16'h012F;    16'd20043: out <= 16'h0683;
    16'd20044: out <= 16'h06D1;    16'd20045: out <= 16'h0A11;    16'd20046: out <= 16'h047F;    16'd20047: out <= 16'h01E4;
    16'd20048: out <= 16'h0423;    16'd20049: out <= 16'h0077;    16'd20050: out <= 16'hFCDC;    16'd20051: out <= 16'h0473;
    16'd20052: out <= 16'h05E5;    16'd20053: out <= 16'h00A4;    16'd20054: out <= 16'h0DB0;    16'd20055: out <= 16'h020E;
    16'd20056: out <= 16'h0941;    16'd20057: out <= 16'h0042;    16'd20058: out <= 16'h07DD;    16'd20059: out <= 16'h0609;
    16'd20060: out <= 16'h045C;    16'd20061: out <= 16'h012B;    16'd20062: out <= 16'hFFF1;    16'd20063: out <= 16'h08FE;
    16'd20064: out <= 16'h0397;    16'd20065: out <= 16'h07FD;    16'd20066: out <= 16'hFEA0;    16'd20067: out <= 16'h0C40;
    16'd20068: out <= 16'h04E8;    16'd20069: out <= 16'h08D7;    16'd20070: out <= 16'h0442;    16'd20071: out <= 16'h00EE;
    16'd20072: out <= 16'hFCDF;    16'd20073: out <= 16'h0450;    16'd20074: out <= 16'h0E65;    16'd20075: out <= 16'hFDE3;
    16'd20076: out <= 16'h02F7;    16'd20077: out <= 16'h0315;    16'd20078: out <= 16'h0544;    16'd20079: out <= 16'h03CD;
    16'd20080: out <= 16'h055A;    16'd20081: out <= 16'h058C;    16'd20082: out <= 16'h0325;    16'd20083: out <= 16'h058B;
    16'd20084: out <= 16'h0419;    16'd20085: out <= 16'h0426;    16'd20086: out <= 16'hFD0F;    16'd20087: out <= 16'h0352;
    16'd20088: out <= 16'h07EC;    16'd20089: out <= 16'h0356;    16'd20090: out <= 16'h0744;    16'd20091: out <= 16'h0229;
    16'd20092: out <= 16'hF6FB;    16'd20093: out <= 16'h0821;    16'd20094: out <= 16'h07F9;    16'd20095: out <= 16'h035F;
    16'd20096: out <= 16'h073F;    16'd20097: out <= 16'h0162;    16'd20098: out <= 16'hFEC5;    16'd20099: out <= 16'h05C6;
    16'd20100: out <= 16'hFE84;    16'd20101: out <= 16'h0A2C;    16'd20102: out <= 16'h0260;    16'd20103: out <= 16'h0A71;
    16'd20104: out <= 16'h09EC;    16'd20105: out <= 16'h07B5;    16'd20106: out <= 16'h04A1;    16'd20107: out <= 16'h0170;
    16'd20108: out <= 16'h0278;    16'd20109: out <= 16'h03DE;    16'd20110: out <= 16'hFF5B;    16'd20111: out <= 16'h05E1;
    16'd20112: out <= 16'h041D;    16'd20113: out <= 16'hFD8A;    16'd20114: out <= 16'h06E1;    16'd20115: out <= 16'h07C1;
    16'd20116: out <= 16'hFC78;    16'd20117: out <= 16'hFE76;    16'd20118: out <= 16'h0051;    16'd20119: out <= 16'h045E;
    16'd20120: out <= 16'hFD37;    16'd20121: out <= 16'h0479;    16'd20122: out <= 16'hFF1E;    16'd20123: out <= 16'h09B6;
    16'd20124: out <= 16'h020E;    16'd20125: out <= 16'hFF99;    16'd20126: out <= 16'h0313;    16'd20127: out <= 16'h03E1;
    16'd20128: out <= 16'h0173;    16'd20129: out <= 16'h0611;    16'd20130: out <= 16'hFFDA;    16'd20131: out <= 16'h011B;
    16'd20132: out <= 16'h08D9;    16'd20133: out <= 16'hFFCA;    16'd20134: out <= 16'h0748;    16'd20135: out <= 16'h03BD;
    16'd20136: out <= 16'hFFF7;    16'd20137: out <= 16'h01D8;    16'd20138: out <= 16'h0261;    16'd20139: out <= 16'h05BC;
    16'd20140: out <= 16'h021F;    16'd20141: out <= 16'h0426;    16'd20142: out <= 16'h0857;    16'd20143: out <= 16'h0D5C;
    16'd20144: out <= 16'hFD0B;    16'd20145: out <= 16'h04B2;    16'd20146: out <= 16'h02E5;    16'd20147: out <= 16'h02EA;
    16'd20148: out <= 16'h092B;    16'd20149: out <= 16'h06B3;    16'd20150: out <= 16'h022D;    16'd20151: out <= 16'h0032;
    16'd20152: out <= 16'h0885;    16'd20153: out <= 16'h0055;    16'd20154: out <= 16'h01B9;    16'd20155: out <= 16'h08D9;
    16'd20156: out <= 16'h04E4;    16'd20157: out <= 16'h031D;    16'd20158: out <= 16'h0228;    16'd20159: out <= 16'h074F;
    16'd20160: out <= 16'hFE84;    16'd20161: out <= 16'h0613;    16'd20162: out <= 16'h0403;    16'd20163: out <= 16'h0296;
    16'd20164: out <= 16'h02BE;    16'd20165: out <= 16'hFCD0;    16'd20166: out <= 16'h04B8;    16'd20167: out <= 16'h05E4;
    16'd20168: out <= 16'h0891;    16'd20169: out <= 16'h062C;    16'd20170: out <= 16'h062F;    16'd20171: out <= 16'h049E;
    16'd20172: out <= 16'h0A6A;    16'd20173: out <= 16'h054B;    16'd20174: out <= 16'h0031;    16'd20175: out <= 16'hFD68;
    16'd20176: out <= 16'h07C0;    16'd20177: out <= 16'h0615;    16'd20178: out <= 16'h02A6;    16'd20179: out <= 16'h01B4;
    16'd20180: out <= 16'hFBAC;    16'd20181: out <= 16'h0806;    16'd20182: out <= 16'h0604;    16'd20183: out <= 16'h0294;
    16'd20184: out <= 16'h0170;    16'd20185: out <= 16'h044A;    16'd20186: out <= 16'h01D1;    16'd20187: out <= 16'h00D3;
    16'd20188: out <= 16'hFC0D;    16'd20189: out <= 16'hF788;    16'd20190: out <= 16'hFBAB;    16'd20191: out <= 16'hFD02;
    16'd20192: out <= 16'hFA1A;    16'd20193: out <= 16'h04A3;    16'd20194: out <= 16'h0158;    16'd20195: out <= 16'h0571;
    16'd20196: out <= 16'h0073;    16'd20197: out <= 16'h05DE;    16'd20198: out <= 16'hFD54;    16'd20199: out <= 16'h01EB;
    16'd20200: out <= 16'h0233;    16'd20201: out <= 16'hFECE;    16'd20202: out <= 16'h00A6;    16'd20203: out <= 16'h0221;
    16'd20204: out <= 16'hF7E0;    16'd20205: out <= 16'h01D5;    16'd20206: out <= 16'h055B;    16'd20207: out <= 16'h075C;
    16'd20208: out <= 16'hFDC1;    16'd20209: out <= 16'hFDA9;    16'd20210: out <= 16'h0235;    16'd20211: out <= 16'hFCE5;
    16'd20212: out <= 16'h0121;    16'd20213: out <= 16'hFF1F;    16'd20214: out <= 16'h00BD;    16'd20215: out <= 16'hF9FB;
    16'd20216: out <= 16'h0606;    16'd20217: out <= 16'hFFE3;    16'd20218: out <= 16'h017C;    16'd20219: out <= 16'h01AE;
    16'd20220: out <= 16'h03B9;    16'd20221: out <= 16'hFAD0;    16'd20222: out <= 16'h032B;    16'd20223: out <= 16'hFD89;
    16'd20224: out <= 16'h039F;    16'd20225: out <= 16'h01F4;    16'd20226: out <= 16'h0B4C;    16'd20227: out <= 16'h0242;
    16'd20228: out <= 16'h03DF;    16'd20229: out <= 16'h0083;    16'd20230: out <= 16'h024F;    16'd20231: out <= 16'h0353;
    16'd20232: out <= 16'hFF2B;    16'd20233: out <= 16'hFC7A;    16'd20234: out <= 16'hFB70;    16'd20235: out <= 16'h020A;
    16'd20236: out <= 16'h0285;    16'd20237: out <= 16'h06C9;    16'd20238: out <= 16'hFF2A;    16'd20239: out <= 16'h00E0;
    16'd20240: out <= 16'h02F6;    16'd20241: out <= 16'hFE15;    16'd20242: out <= 16'h0354;    16'd20243: out <= 16'hFFCF;
    16'd20244: out <= 16'hFDA1;    16'd20245: out <= 16'hFE51;    16'd20246: out <= 16'h00A4;    16'd20247: out <= 16'hFE7A;
    16'd20248: out <= 16'hF83D;    16'd20249: out <= 16'hFF9F;    16'd20250: out <= 16'hFD71;    16'd20251: out <= 16'h053B;
    16'd20252: out <= 16'h04DA;    16'd20253: out <= 16'h02D7;    16'd20254: out <= 16'hFF5B;    16'd20255: out <= 16'h0570;
    16'd20256: out <= 16'h01BE;    16'd20257: out <= 16'h071B;    16'd20258: out <= 16'h0859;    16'd20259: out <= 16'h0376;
    16'd20260: out <= 16'h001A;    16'd20261: out <= 16'h08A9;    16'd20262: out <= 16'hFCB2;    16'd20263: out <= 16'h043D;
    16'd20264: out <= 16'h003B;    16'd20265: out <= 16'h0268;    16'd20266: out <= 16'h06AB;    16'd20267: out <= 16'h0822;
    16'd20268: out <= 16'h05BB;    16'd20269: out <= 16'h04F4;    16'd20270: out <= 16'h01C0;    16'd20271: out <= 16'h03D3;
    16'd20272: out <= 16'h04F6;    16'd20273: out <= 16'h0016;    16'd20274: out <= 16'h05CE;    16'd20275: out <= 16'hFF56;
    16'd20276: out <= 16'h017D;    16'd20277: out <= 16'h060C;    16'd20278: out <= 16'h041F;    16'd20279: out <= 16'h005E;
    16'd20280: out <= 16'h063E;    16'd20281: out <= 16'h023E;    16'd20282: out <= 16'h00DE;    16'd20283: out <= 16'hFEAD;
    16'd20284: out <= 16'h0717;    16'd20285: out <= 16'h0972;    16'd20286: out <= 16'h062B;    16'd20287: out <= 16'h0099;
    16'd20288: out <= 16'h02F5;    16'd20289: out <= 16'hFC3B;    16'd20290: out <= 16'h026E;    16'd20291: out <= 16'h09F3;
    16'd20292: out <= 16'h0281;    16'd20293: out <= 16'h02BA;    16'd20294: out <= 16'hFC75;    16'd20295: out <= 16'hFD49;
    16'd20296: out <= 16'h0519;    16'd20297: out <= 16'hFDC8;    16'd20298: out <= 16'h0469;    16'd20299: out <= 16'h06D5;
    16'd20300: out <= 16'h02B6;    16'd20301: out <= 16'h0839;    16'd20302: out <= 16'hFBB7;    16'd20303: out <= 16'h01D9;
    16'd20304: out <= 16'h052C;    16'd20305: out <= 16'hFBFB;    16'd20306: out <= 16'hF9D5;    16'd20307: out <= 16'h0436;
    16'd20308: out <= 16'h04F7;    16'd20309: out <= 16'h0148;    16'd20310: out <= 16'hFFBA;    16'd20311: out <= 16'h0009;
    16'd20312: out <= 16'h0955;    16'd20313: out <= 16'h0539;    16'd20314: out <= 16'h06D8;    16'd20315: out <= 16'h02C8;
    16'd20316: out <= 16'h04B6;    16'd20317: out <= 16'h059B;    16'd20318: out <= 16'h04BC;    16'd20319: out <= 16'h02C0;
    16'd20320: out <= 16'h0540;    16'd20321: out <= 16'h0583;    16'd20322: out <= 16'hFB77;    16'd20323: out <= 16'h02C6;
    16'd20324: out <= 16'h04A9;    16'd20325: out <= 16'h0442;    16'd20326: out <= 16'h0562;    16'd20327: out <= 16'h059B;
    16'd20328: out <= 16'h0BD0;    16'd20329: out <= 16'h0279;    16'd20330: out <= 16'h0278;    16'd20331: out <= 16'h060E;
    16'd20332: out <= 16'h07E8;    16'd20333: out <= 16'h0225;    16'd20334: out <= 16'hFAD1;    16'd20335: out <= 16'h05B4;
    16'd20336: out <= 16'h073B;    16'd20337: out <= 16'h03EB;    16'd20338: out <= 16'h0524;    16'd20339: out <= 16'h066B;
    16'd20340: out <= 16'h0977;    16'd20341: out <= 16'h0383;    16'd20342: out <= 16'h0219;    16'd20343: out <= 16'h0484;
    16'd20344: out <= 16'h0724;    16'd20345: out <= 16'h069B;    16'd20346: out <= 16'h062C;    16'd20347: out <= 16'hFDDA;
    16'd20348: out <= 16'h00F9;    16'd20349: out <= 16'h0432;    16'd20350: out <= 16'h03C6;    16'd20351: out <= 16'h0A4B;
    16'd20352: out <= 16'h00B7;    16'd20353: out <= 16'h02E8;    16'd20354: out <= 16'h013F;    16'd20355: out <= 16'h09D6;
    16'd20356: out <= 16'h04A8;    16'd20357: out <= 16'h01C8;    16'd20358: out <= 16'hFE65;    16'd20359: out <= 16'h0292;
    16'd20360: out <= 16'h018F;    16'd20361: out <= 16'h020B;    16'd20362: out <= 16'h01C1;    16'd20363: out <= 16'h001C;
    16'd20364: out <= 16'h0374;    16'd20365: out <= 16'h02F3;    16'd20366: out <= 16'h0045;    16'd20367: out <= 16'h021C;
    16'd20368: out <= 16'h0439;    16'd20369: out <= 16'h02E3;    16'd20370: out <= 16'h0604;    16'd20371: out <= 16'h029C;
    16'd20372: out <= 16'h0385;    16'd20373: out <= 16'hFFC1;    16'd20374: out <= 16'h04DD;    16'd20375: out <= 16'h0281;
    16'd20376: out <= 16'h05EA;    16'd20377: out <= 16'h00C6;    16'd20378: out <= 16'h05E3;    16'd20379: out <= 16'h09D9;
    16'd20380: out <= 16'h050E;    16'd20381: out <= 16'h0592;    16'd20382: out <= 16'h09DD;    16'd20383: out <= 16'h0A39;
    16'd20384: out <= 16'h0AE6;    16'd20385: out <= 16'h071B;    16'd20386: out <= 16'h0319;    16'd20387: out <= 16'hFF7D;
    16'd20388: out <= 16'h00AD;    16'd20389: out <= 16'h029A;    16'd20390: out <= 16'h03C4;    16'd20391: out <= 16'hFFFE;
    16'd20392: out <= 16'h0C21;    16'd20393: out <= 16'hFE24;    16'd20394: out <= 16'h0843;    16'd20395: out <= 16'hFEB6;
    16'd20396: out <= 16'h0356;    16'd20397: out <= 16'h067C;    16'd20398: out <= 16'h06A8;    16'd20399: out <= 16'hFAE6;
    16'd20400: out <= 16'h048C;    16'd20401: out <= 16'h0C34;    16'd20402: out <= 16'h0385;    16'd20403: out <= 16'hFA4C;
    16'd20404: out <= 16'h0329;    16'd20405: out <= 16'hFE37;    16'd20406: out <= 16'h04D5;    16'd20407: out <= 16'h0483;
    16'd20408: out <= 16'h083E;    16'd20409: out <= 16'h0838;    16'd20410: out <= 16'h0324;    16'd20411: out <= 16'h0B37;
    16'd20412: out <= 16'h01C7;    16'd20413: out <= 16'hFEC4;    16'd20414: out <= 16'h075B;    16'd20415: out <= 16'h048F;
    16'd20416: out <= 16'h05A9;    16'd20417: out <= 16'h0068;    16'd20418: out <= 16'h0603;    16'd20419: out <= 16'h02C8;
    16'd20420: out <= 16'h0B6E;    16'd20421: out <= 16'h07F9;    16'd20422: out <= 16'h041E;    16'd20423: out <= 16'h03E1;
    16'd20424: out <= 16'hFF16;    16'd20425: out <= 16'h0663;    16'd20426: out <= 16'hFE84;    16'd20427: out <= 16'hFE00;
    16'd20428: out <= 16'h0086;    16'd20429: out <= 16'h03A0;    16'd20430: out <= 16'h0186;    16'd20431: out <= 16'h0554;
    16'd20432: out <= 16'h04D1;    16'd20433: out <= 16'hFF68;    16'd20434: out <= 16'h0439;    16'd20435: out <= 16'h057B;
    16'd20436: out <= 16'h05FA;    16'd20437: out <= 16'h02CF;    16'd20438: out <= 16'h0165;    16'd20439: out <= 16'h0168;
    16'd20440: out <= 16'h00E5;    16'd20441: out <= 16'h02B3;    16'd20442: out <= 16'hFE3F;    16'd20443: out <= 16'h003F;
    16'd20444: out <= 16'h0522;    16'd20445: out <= 16'hFF35;    16'd20446: out <= 16'hFEB8;    16'd20447: out <= 16'hFD31;
    16'd20448: out <= 16'h034A;    16'd20449: out <= 16'hFD87;    16'd20450: out <= 16'hFD8B;    16'd20451: out <= 16'h0217;
    16'd20452: out <= 16'h0215;    16'd20453: out <= 16'hFCCE;    16'd20454: out <= 16'hFDD9;    16'd20455: out <= 16'hFD59;
    16'd20456: out <= 16'h0681;    16'd20457: out <= 16'hFBB7;    16'd20458: out <= 16'h003C;    16'd20459: out <= 16'h0755;
    16'd20460: out <= 16'h0239;    16'd20461: out <= 16'h067A;    16'd20462: out <= 16'hFE38;    16'd20463: out <= 16'h01CA;
    16'd20464: out <= 16'h001A;    16'd20465: out <= 16'hFD4E;    16'd20466: out <= 16'h006B;    16'd20467: out <= 16'hFEF8;
    16'd20468: out <= 16'h0587;    16'd20469: out <= 16'hFE9F;    16'd20470: out <= 16'h001D;    16'd20471: out <= 16'hFCF7;
    16'd20472: out <= 16'hFB4D;    16'd20473: out <= 16'h0517;    16'd20474: out <= 16'hFCA7;    16'd20475: out <= 16'hFF11;
    16'd20476: out <= 16'h06A2;    16'd20477: out <= 16'h022E;    16'd20478: out <= 16'hFC5B;    16'd20479: out <= 16'hF97B;
    16'd20480: out <= 16'hFF59;    16'd20481: out <= 16'h03A0;    16'd20482: out <= 16'h0438;    16'd20483: out <= 16'hFAEC;
    16'd20484: out <= 16'h0027;    16'd20485: out <= 16'h004C;    16'd20486: out <= 16'h00D4;    16'd20487: out <= 16'h0151;
    16'd20488: out <= 16'h00B3;    16'd20489: out <= 16'hFA63;    16'd20490: out <= 16'hFE70;    16'd20491: out <= 16'hFEBF;
    16'd20492: out <= 16'h03E5;    16'd20493: out <= 16'hFF9C;    16'd20494: out <= 16'h00CF;    16'd20495: out <= 16'hFEEA;
    16'd20496: out <= 16'h066C;    16'd20497: out <= 16'h0320;    16'd20498: out <= 16'h04EF;    16'd20499: out <= 16'h02F9;
    16'd20500: out <= 16'h02CB;    16'd20501: out <= 16'h01AA;    16'd20502: out <= 16'hFD2A;    16'd20503: out <= 16'h0000;
    16'd20504: out <= 16'hFFC2;    16'd20505: out <= 16'hFD40;    16'd20506: out <= 16'h09A4;    16'd20507: out <= 16'h02CA;
    16'd20508: out <= 16'h004B;    16'd20509: out <= 16'h022C;    16'd20510: out <= 16'h048A;    16'd20511: out <= 16'h01A0;
    16'd20512: out <= 16'hFDA3;    16'd20513: out <= 16'h04BA;    16'd20514: out <= 16'h0DE2;    16'd20515: out <= 16'h06A0;
    16'd20516: out <= 16'hFF28;    16'd20517: out <= 16'h0540;    16'd20518: out <= 16'h05E0;    16'd20519: out <= 16'hFE98;
    16'd20520: out <= 16'h027B;    16'd20521: out <= 16'h0118;    16'd20522: out <= 16'h0649;    16'd20523: out <= 16'h0639;
    16'd20524: out <= 16'h07BA;    16'd20525: out <= 16'h086C;    16'd20526: out <= 16'h0907;    16'd20527: out <= 16'h0311;
    16'd20528: out <= 16'h04D4;    16'd20529: out <= 16'h00A4;    16'd20530: out <= 16'hFEF6;    16'd20531: out <= 16'h03DD;
    16'd20532: out <= 16'hFF8F;    16'd20533: out <= 16'h0629;    16'd20534: out <= 16'h08C2;    16'd20535: out <= 16'hF744;
    16'd20536: out <= 16'h09F1;    16'd20537: out <= 16'h03CE;    16'd20538: out <= 16'h0A8C;    16'd20539: out <= 16'h0330;
    16'd20540: out <= 16'h099E;    16'd20541: out <= 16'h069B;    16'd20542: out <= 16'h05DC;    16'd20543: out <= 16'hFD7D;
    16'd20544: out <= 16'h033C;    16'd20545: out <= 16'h013E;    16'd20546: out <= 16'h057B;    16'd20547: out <= 16'h03D3;
    16'd20548: out <= 16'h029E;    16'd20549: out <= 16'h02DE;    16'd20550: out <= 16'hFD34;    16'd20551: out <= 16'h02B3;
    16'd20552: out <= 16'h09B3;    16'd20553: out <= 16'h0353;    16'd20554: out <= 16'h08E8;    16'd20555: out <= 16'h0187;
    16'd20556: out <= 16'h0693;    16'd20557: out <= 16'h011C;    16'd20558: out <= 16'hFC48;    16'd20559: out <= 16'h0106;
    16'd20560: out <= 16'h05B1;    16'd20561: out <= 16'h0160;    16'd20562: out <= 16'h0388;    16'd20563: out <= 16'h0837;
    16'd20564: out <= 16'h01A9;    16'd20565: out <= 16'h0534;    16'd20566: out <= 16'h095B;    16'd20567: out <= 16'h0978;
    16'd20568: out <= 16'h075F;    16'd20569: out <= 16'h0555;    16'd20570: out <= 16'h01EB;    16'd20571: out <= 16'h036C;
    16'd20572: out <= 16'hFCD8;    16'd20573: out <= 16'h03CF;    16'd20574: out <= 16'h01EA;    16'd20575: out <= 16'h0159;
    16'd20576: out <= 16'hF910;    16'd20577: out <= 16'h033B;    16'd20578: out <= 16'h030E;    16'd20579: out <= 16'h0A97;
    16'd20580: out <= 16'hF6D5;    16'd20581: out <= 16'h000D;    16'd20582: out <= 16'h086B;    16'd20583: out <= 16'h0258;
    16'd20584: out <= 16'h009D;    16'd20585: out <= 16'h09B3;    16'd20586: out <= 16'h02FC;    16'd20587: out <= 16'h08BB;
    16'd20588: out <= 16'h05B7;    16'd20589: out <= 16'h0825;    16'd20590: out <= 16'h0051;    16'd20591: out <= 16'h0829;
    16'd20592: out <= 16'hFCEE;    16'd20593: out <= 16'h0032;    16'd20594: out <= 16'h018D;    16'd20595: out <= 16'h0436;
    16'd20596: out <= 16'h0225;    16'd20597: out <= 16'h0356;    16'd20598: out <= 16'h05A5;    16'd20599: out <= 16'h0721;
    16'd20600: out <= 16'h0102;    16'd20601: out <= 16'h074B;    16'd20602: out <= 16'h029B;    16'd20603: out <= 16'h0001;
    16'd20604: out <= 16'h02FC;    16'd20605: out <= 16'h04FF;    16'd20606: out <= 16'h0388;    16'd20607: out <= 16'h0715;
    16'd20608: out <= 16'h0992;    16'd20609: out <= 16'h060C;    16'd20610: out <= 16'hFF0D;    16'd20611: out <= 16'h00A4;
    16'd20612: out <= 16'h023A;    16'd20613: out <= 16'h0499;    16'd20614: out <= 16'h0C41;    16'd20615: out <= 16'h0763;
    16'd20616: out <= 16'h0C75;    16'd20617: out <= 16'hFD8D;    16'd20618: out <= 16'h0326;    16'd20619: out <= 16'h034E;
    16'd20620: out <= 16'h0146;    16'd20621: out <= 16'h0639;    16'd20622: out <= 16'h0579;    16'd20623: out <= 16'h037F;
    16'd20624: out <= 16'h0A4C;    16'd20625: out <= 16'h056C;    16'd20626: out <= 16'h0175;    16'd20627: out <= 16'h03A2;
    16'd20628: out <= 16'h0602;    16'd20629: out <= 16'h009A;    16'd20630: out <= 16'h067F;    16'd20631: out <= 16'h0284;
    16'd20632: out <= 16'h01ED;    16'd20633: out <= 16'h0415;    16'd20634: out <= 16'h03DD;    16'd20635: out <= 16'h02ED;
    16'd20636: out <= 16'h0383;    16'd20637: out <= 16'hFCEB;    16'd20638: out <= 16'hFB61;    16'd20639: out <= 16'h05AA;
    16'd20640: out <= 16'h01EF;    16'd20641: out <= 16'h04DC;    16'd20642: out <= 16'h0676;    16'd20643: out <= 16'hF432;
    16'd20644: out <= 16'h04E0;    16'd20645: out <= 16'hFE15;    16'd20646: out <= 16'h08C7;    16'd20647: out <= 16'h09DC;
    16'd20648: out <= 16'h0790;    16'd20649: out <= 16'h0DC7;    16'd20650: out <= 16'h0557;    16'd20651: out <= 16'h0AE4;
    16'd20652: out <= 16'h0008;    16'd20653: out <= 16'h085B;    16'd20654: out <= 16'h0AAE;    16'd20655: out <= 16'h069B;
    16'd20656: out <= 16'h0369;    16'd20657: out <= 16'h0402;    16'd20658: out <= 16'h08C8;    16'd20659: out <= 16'hF961;
    16'd20660: out <= 16'h0794;    16'd20661: out <= 16'h05FB;    16'd20662: out <= 16'h073E;    16'd20663: out <= 16'h017D;
    16'd20664: out <= 16'h06A5;    16'd20665: out <= 16'h057B;    16'd20666: out <= 16'h0290;    16'd20667: out <= 16'hFF57;
    16'd20668: out <= 16'h015E;    16'd20669: out <= 16'h0716;    16'd20670: out <= 16'h0597;    16'd20671: out <= 16'h034B;
    16'd20672: out <= 16'h0379;    16'd20673: out <= 16'h0909;    16'd20674: out <= 16'h00CD;    16'd20675: out <= 16'h0149;
    16'd20676: out <= 16'h052D;    16'd20677: out <= 16'h05E8;    16'd20678: out <= 16'h0A97;    16'd20679: out <= 16'h05D9;
    16'd20680: out <= 16'hFF80;    16'd20681: out <= 16'h0396;    16'd20682: out <= 16'h0300;    16'd20683: out <= 16'h02A0;
    16'd20684: out <= 16'h0639;    16'd20685: out <= 16'h0430;    16'd20686: out <= 16'hFE0F;    16'd20687: out <= 16'h0C1E;
    16'd20688: out <= 16'h07D9;    16'd20689: out <= 16'hFA4D;    16'd20690: out <= 16'h056C;    16'd20691: out <= 16'h0743;
    16'd20692: out <= 16'h02A8;    16'd20693: out <= 16'h0301;    16'd20694: out <= 16'h0054;    16'd20695: out <= 16'hFF1E;
    16'd20696: out <= 16'h040F;    16'd20697: out <= 16'h0125;    16'd20698: out <= 16'h015F;    16'd20699: out <= 16'h0602;
    16'd20700: out <= 16'hFF33;    16'd20701: out <= 16'hFF29;    16'd20702: out <= 16'h0029;    16'd20703: out <= 16'hFDA4;
    16'd20704: out <= 16'h01B8;    16'd20705: out <= 16'h03C5;    16'd20706: out <= 16'hFF38;    16'd20707: out <= 16'h00AC;
    16'd20708: out <= 16'hFB6D;    16'd20709: out <= 16'h012C;    16'd20710: out <= 16'h000D;    16'd20711: out <= 16'hFA9C;
    16'd20712: out <= 16'h011A;    16'd20713: out <= 16'h0002;    16'd20714: out <= 16'h004D;    16'd20715: out <= 16'hFB32;
    16'd20716: out <= 16'hFCA9;    16'd20717: out <= 16'hFDAC;    16'd20718: out <= 16'h0556;    16'd20719: out <= 16'h05BB;
    16'd20720: out <= 16'hFDC6;    16'd20721: out <= 16'h0291;    16'd20722: out <= 16'h01EB;    16'd20723: out <= 16'hFEB6;
    16'd20724: out <= 16'hFDE3;    16'd20725: out <= 16'hFFC7;    16'd20726: out <= 16'hFFCE;    16'd20727: out <= 16'h0086;
    16'd20728: out <= 16'hF98A;    16'd20729: out <= 16'hFF16;    16'd20730: out <= 16'h0095;    16'd20731: out <= 16'hFA58;
    16'd20732: out <= 16'h03A0;    16'd20733: out <= 16'h0062;    16'd20734: out <= 16'h0299;    16'd20735: out <= 16'hF65C;
    16'd20736: out <= 16'hF844;    16'd20737: out <= 16'hFD3B;    16'd20738: out <= 16'hFDD9;    16'd20739: out <= 16'hFDF7;
    16'd20740: out <= 16'hFFBE;    16'd20741: out <= 16'hFC1F;    16'd20742: out <= 16'h0731;    16'd20743: out <= 16'hF935;
    16'd20744: out <= 16'h000C;    16'd20745: out <= 16'hFF5A;    16'd20746: out <= 16'h058B;    16'd20747: out <= 16'h010C;
    16'd20748: out <= 16'hF66A;    16'd20749: out <= 16'h0563;    16'd20750: out <= 16'hFFCF;    16'd20751: out <= 16'hFBEB;
    16'd20752: out <= 16'h03DA;    16'd20753: out <= 16'hFBF6;    16'd20754: out <= 16'hFCAE;    16'd20755: out <= 16'h01BC;
    16'd20756: out <= 16'hFEB2;    16'd20757: out <= 16'hF717;    16'd20758: out <= 16'hFE10;    16'd20759: out <= 16'h020D;
    16'd20760: out <= 16'hF726;    16'd20761: out <= 16'h09EC;    16'd20762: out <= 16'h009B;    16'd20763: out <= 16'h0979;
    16'd20764: out <= 16'hFE5E;    16'd20765: out <= 16'h046D;    16'd20766: out <= 16'hFF86;    16'd20767: out <= 16'hFF27;
    16'd20768: out <= 16'hFEEB;    16'd20769: out <= 16'h0609;    16'd20770: out <= 16'h0904;    16'd20771: out <= 16'h0677;
    16'd20772: out <= 16'h052F;    16'd20773: out <= 16'h040B;    16'd20774: out <= 16'h0A8F;    16'd20775: out <= 16'h0308;
    16'd20776: out <= 16'h0A91;    16'd20777: out <= 16'h02AC;    16'd20778: out <= 16'hFDF2;    16'd20779: out <= 16'h009B;
    16'd20780: out <= 16'h0216;    16'd20781: out <= 16'h0254;    16'd20782: out <= 16'h0524;    16'd20783: out <= 16'h0904;
    16'd20784: out <= 16'h034E;    16'd20785: out <= 16'hFFEE;    16'd20786: out <= 16'h0115;    16'd20787: out <= 16'h0675;
    16'd20788: out <= 16'h015F;    16'd20789: out <= 16'hFD55;    16'd20790: out <= 16'h01EC;    16'd20791: out <= 16'h0BE7;
    16'd20792: out <= 16'h0870;    16'd20793: out <= 16'h0268;    16'd20794: out <= 16'h0915;    16'd20795: out <= 16'h03DA;
    16'd20796: out <= 16'hFF85;    16'd20797: out <= 16'hFF7A;    16'd20798: out <= 16'h00D0;    16'd20799: out <= 16'h06B5;
    16'd20800: out <= 16'h0D49;    16'd20801: out <= 16'hFD50;    16'd20802: out <= 16'h07C5;    16'd20803: out <= 16'h0405;
    16'd20804: out <= 16'h0523;    16'd20805: out <= 16'h02D3;    16'd20806: out <= 16'h06B6;    16'd20807: out <= 16'h02EB;
    16'd20808: out <= 16'h030D;    16'd20809: out <= 16'h0CCB;    16'd20810: out <= 16'h07F4;    16'd20811: out <= 16'h0970;
    16'd20812: out <= 16'h000C;    16'd20813: out <= 16'hFBD6;    16'd20814: out <= 16'hFBAB;    16'd20815: out <= 16'h005C;
    16'd20816: out <= 16'h0843;    16'd20817: out <= 16'h0138;    16'd20818: out <= 16'h03E6;    16'd20819: out <= 16'h069E;
    16'd20820: out <= 16'h03DD;    16'd20821: out <= 16'h0477;    16'd20822: out <= 16'h08AF;    16'd20823: out <= 16'h05B1;
    16'd20824: out <= 16'h00A5;    16'd20825: out <= 16'h088C;    16'd20826: out <= 16'h069C;    16'd20827: out <= 16'h05F5;
    16'd20828: out <= 16'h01CD;    16'd20829: out <= 16'hFFC1;    16'd20830: out <= 16'h0205;    16'd20831: out <= 16'h08E5;
    16'd20832: out <= 16'h0281;    16'd20833: out <= 16'h0591;    16'd20834: out <= 16'h0378;    16'd20835: out <= 16'hFFAC;
    16'd20836: out <= 16'hFC28;    16'd20837: out <= 16'h0021;    16'd20838: out <= 16'h03C9;    16'd20839: out <= 16'h08D1;
    16'd20840: out <= 16'h0068;    16'd20841: out <= 16'h07FA;    16'd20842: out <= 16'h0511;    16'd20843: out <= 16'h02E8;
    16'd20844: out <= 16'hFBFB;    16'd20845: out <= 16'hFA90;    16'd20846: out <= 16'h0768;    16'd20847: out <= 16'h0649;
    16'd20848: out <= 16'h02D2;    16'd20849: out <= 16'h0772;    16'd20850: out <= 16'h029F;    16'd20851: out <= 16'h06A6;
    16'd20852: out <= 16'h008C;    16'd20853: out <= 16'hFC59;    16'd20854: out <= 16'h0380;    16'd20855: out <= 16'h051E;
    16'd20856: out <= 16'h0647;    16'd20857: out <= 16'h097A;    16'd20858: out <= 16'h0521;    16'd20859: out <= 16'h0383;
    16'd20860: out <= 16'h06E5;    16'd20861: out <= 16'hFE69;    16'd20862: out <= 16'h0704;    16'd20863: out <= 16'h063D;
    16'd20864: out <= 16'h085F;    16'd20865: out <= 16'h0138;    16'd20866: out <= 16'h01DA;    16'd20867: out <= 16'h0490;
    16'd20868: out <= 16'hFD4D;    16'd20869: out <= 16'h0646;    16'd20870: out <= 16'h0210;    16'd20871: out <= 16'h00D5;
    16'd20872: out <= 16'h012C;    16'd20873: out <= 16'h01D8;    16'd20874: out <= 16'h000D;    16'd20875: out <= 16'hFE71;
    16'd20876: out <= 16'h0458;    16'd20877: out <= 16'h027D;    16'd20878: out <= 16'h0152;    16'd20879: out <= 16'h000F;
    16'd20880: out <= 16'h0429;    16'd20881: out <= 16'h0533;    16'd20882: out <= 16'h0905;    16'd20883: out <= 16'h047F;
    16'd20884: out <= 16'h06C7;    16'd20885: out <= 16'h09A2;    16'd20886: out <= 16'hFDCA;    16'd20887: out <= 16'h0151;
    16'd20888: out <= 16'h0278;    16'd20889: out <= 16'h0001;    16'd20890: out <= 16'h0B0C;    16'd20891: out <= 16'h095E;
    16'd20892: out <= 16'hFF98;    16'd20893: out <= 16'h0B38;    16'd20894: out <= 16'h0862;    16'd20895: out <= 16'h03D6;
    16'd20896: out <= 16'h0566;    16'd20897: out <= 16'h01F2;    16'd20898: out <= 16'hFF0E;    16'd20899: out <= 16'hFD4C;
    16'd20900: out <= 16'h076D;    16'd20901: out <= 16'h09E5;    16'd20902: out <= 16'h0105;    16'd20903: out <= 16'hFF65;
    16'd20904: out <= 16'h0649;    16'd20905: out <= 16'h06E9;    16'd20906: out <= 16'h000E;    16'd20907: out <= 16'h033B;
    16'd20908: out <= 16'h02A4;    16'd20909: out <= 16'h02CD;    16'd20910: out <= 16'h0237;    16'd20911: out <= 16'h02AF;
    16'd20912: out <= 16'h024E;    16'd20913: out <= 16'h0BAE;    16'd20914: out <= 16'hFF92;    16'd20915: out <= 16'h011D;
    16'd20916: out <= 16'h04C4;    16'd20917: out <= 16'h02FC;    16'd20918: out <= 16'h0796;    16'd20919: out <= 16'h0710;
    16'd20920: out <= 16'h02AB;    16'd20921: out <= 16'h03E1;    16'd20922: out <= 16'h01F1;    16'd20923: out <= 16'h065D;
    16'd20924: out <= 16'h05B7;    16'd20925: out <= 16'h08FD;    16'd20926: out <= 16'h0450;    16'd20927: out <= 16'h04D8;
    16'd20928: out <= 16'h04F7;    16'd20929: out <= 16'h02C6;    16'd20930: out <= 16'h06D3;    16'd20931: out <= 16'h00A9;
    16'd20932: out <= 16'h032C;    16'd20933: out <= 16'hFEB9;    16'd20934: out <= 16'h0422;    16'd20935: out <= 16'h03DE;
    16'd20936: out <= 16'hFEDD;    16'd20937: out <= 16'h0634;    16'd20938: out <= 16'h0737;    16'd20939: out <= 16'h04F6;
    16'd20940: out <= 16'h000A;    16'd20941: out <= 16'hFD82;    16'd20942: out <= 16'h0997;    16'd20943: out <= 16'h099B;
    16'd20944: out <= 16'h05AA;    16'd20945: out <= 16'h0116;    16'd20946: out <= 16'h0311;    16'd20947: out <= 16'h0640;
    16'd20948: out <= 16'h08FA;    16'd20949: out <= 16'h0A7B;    16'd20950: out <= 16'h05B1;    16'd20951: out <= 16'hFC53;
    16'd20952: out <= 16'h0684;    16'd20953: out <= 16'h04FC;    16'd20954: out <= 16'h01C3;    16'd20955: out <= 16'h0179;
    16'd20956: out <= 16'hFF79;    16'd20957: out <= 16'h0350;    16'd20958: out <= 16'h00BE;    16'd20959: out <= 16'h04E9;
    16'd20960: out <= 16'h0064;    16'd20961: out <= 16'hF580;    16'd20962: out <= 16'hFB7D;    16'd20963: out <= 16'hFE1E;
    16'd20964: out <= 16'h0693;    16'd20965: out <= 16'h01AE;    16'd20966: out <= 16'h0516;    16'd20967: out <= 16'h0479;
    16'd20968: out <= 16'hFD84;    16'd20969: out <= 16'h01FC;    16'd20970: out <= 16'hFEF0;    16'd20971: out <= 16'h0430;
    16'd20972: out <= 16'h028D;    16'd20973: out <= 16'hFAD9;    16'd20974: out <= 16'hFC35;    16'd20975: out <= 16'hFECE;
    16'd20976: out <= 16'h00AF;    16'd20977: out <= 16'h000C;    16'd20978: out <= 16'h04CD;    16'd20979: out <= 16'h089A;
    16'd20980: out <= 16'hFF52;    16'd20981: out <= 16'hFD46;    16'd20982: out <= 16'hFEC1;    16'd20983: out <= 16'hFAEE;
    16'd20984: out <= 16'hF900;    16'd20985: out <= 16'h0529;    16'd20986: out <= 16'h005F;    16'd20987: out <= 16'hFB74;
    16'd20988: out <= 16'hF485;    16'd20989: out <= 16'hFBBA;    16'd20990: out <= 16'hFC82;    16'd20991: out <= 16'hFF3E;
    16'd20992: out <= 16'hFF54;    16'd20993: out <= 16'h00E3;    16'd20994: out <= 16'h03C8;    16'd20995: out <= 16'h05C4;
    16'd20996: out <= 16'h03BE;    16'd20997: out <= 16'h0227;    16'd20998: out <= 16'hFB4F;    16'd20999: out <= 16'h0188;
    16'd21000: out <= 16'hFCFC;    16'd21001: out <= 16'h0168;    16'd21002: out <= 16'h0291;    16'd21003: out <= 16'h0293;
    16'd21004: out <= 16'h042C;    16'd21005: out <= 16'hFB50;    16'd21006: out <= 16'h0366;    16'd21007: out <= 16'h07CE;
    16'd21008: out <= 16'h012F;    16'd21009: out <= 16'h02D2;    16'd21010: out <= 16'h0903;    16'd21011: out <= 16'hFE99;
    16'd21012: out <= 16'h03B2;    16'd21013: out <= 16'hFCA0;    16'd21014: out <= 16'h0171;    16'd21015: out <= 16'hFB21;
    16'd21016: out <= 16'hFEC4;    16'd21017: out <= 16'h0DBF;    16'd21018: out <= 16'h06C6;    16'd21019: out <= 16'hFEBA;
    16'd21020: out <= 16'h000C;    16'd21021: out <= 16'h0641;    16'd21022: out <= 16'h02FA;    16'd21023: out <= 16'h08B6;
    16'd21024: out <= 16'hFCEA;    16'd21025: out <= 16'h0574;    16'd21026: out <= 16'h095C;    16'd21027: out <= 16'h0471;
    16'd21028: out <= 16'hFFD2;    16'd21029: out <= 16'h03C0;    16'd21030: out <= 16'h05E3;    16'd21031: out <= 16'h06F9;
    16'd21032: out <= 16'h09AA;    16'd21033: out <= 16'hFF1A;    16'd21034: out <= 16'h0281;    16'd21035: out <= 16'h0258;
    16'd21036: out <= 16'h0538;    16'd21037: out <= 16'h06C2;    16'd21038: out <= 16'h01E3;    16'd21039: out <= 16'h03D5;
    16'd21040: out <= 16'h0424;    16'd21041: out <= 16'h0F5F;    16'd21042: out <= 16'h01C3;    16'd21043: out <= 16'h018E;
    16'd21044: out <= 16'h051F;    16'd21045: out <= 16'h00DE;    16'd21046: out <= 16'h083C;    16'd21047: out <= 16'h0646;
    16'd21048: out <= 16'h0300;    16'd21049: out <= 16'h037E;    16'd21050: out <= 16'h03BE;    16'd21051: out <= 16'h083F;
    16'd21052: out <= 16'hFFA9;    16'd21053: out <= 16'h0142;    16'd21054: out <= 16'h025C;    16'd21055: out <= 16'hFF3A;
    16'd21056: out <= 16'h0876;    16'd21057: out <= 16'h058F;    16'd21058: out <= 16'h0602;    16'd21059: out <= 16'hF600;
    16'd21060: out <= 16'h04BE;    16'd21061: out <= 16'h03E3;    16'd21062: out <= 16'h02EB;    16'd21063: out <= 16'h03AD;
    16'd21064: out <= 16'h0608;    16'd21065: out <= 16'hFE79;    16'd21066: out <= 16'h09ED;    16'd21067: out <= 16'h08F5;
    16'd21068: out <= 16'hF916;    16'd21069: out <= 16'hFF6F;    16'd21070: out <= 16'hFF4C;    16'd21071: out <= 16'h021A;
    16'd21072: out <= 16'hFF00;    16'd21073: out <= 16'hFA50;    16'd21074: out <= 16'hFCB6;    16'd21075: out <= 16'hFF5F;
    16'd21076: out <= 16'hFDB2;    16'd21077: out <= 16'h03CC;    16'd21078: out <= 16'h0A5A;    16'd21079: out <= 16'h02AA;
    16'd21080: out <= 16'h05B7;    16'd21081: out <= 16'h0615;    16'd21082: out <= 16'h01C1;    16'd21083: out <= 16'h0283;
    16'd21084: out <= 16'h0183;    16'd21085: out <= 16'h0224;    16'd21086: out <= 16'hFFB8;    16'd21087: out <= 16'h01FE;
    16'd21088: out <= 16'h003A;    16'd21089: out <= 16'h02AA;    16'd21090: out <= 16'h0059;    16'd21091: out <= 16'h0492;
    16'd21092: out <= 16'h0783;    16'd21093: out <= 16'h0229;    16'd21094: out <= 16'h02E7;    16'd21095: out <= 16'h04E4;
    16'd21096: out <= 16'hFC9A;    16'd21097: out <= 16'h014A;    16'd21098: out <= 16'h0629;    16'd21099: out <= 16'h07E9;
    16'd21100: out <= 16'h0538;    16'd21101: out <= 16'h070E;    16'd21102: out <= 16'hFA87;    16'd21103: out <= 16'h067D;
    16'd21104: out <= 16'h0966;    16'd21105: out <= 16'h07D9;    16'd21106: out <= 16'h0AB0;    16'd21107: out <= 16'h046D;
    16'd21108: out <= 16'h08C1;    16'd21109: out <= 16'h05AF;    16'd21110: out <= 16'hFF59;    16'd21111: out <= 16'h003B;
    16'd21112: out <= 16'h034A;    16'd21113: out <= 16'hFE95;    16'd21114: out <= 16'h03E1;    16'd21115: out <= 16'hFCF4;
    16'd21116: out <= 16'h0B7A;    16'd21117: out <= 16'h0784;    16'd21118: out <= 16'h0823;    16'd21119: out <= 16'h0941;
    16'd21120: out <= 16'h02DB;    16'd21121: out <= 16'h003D;    16'd21122: out <= 16'h0208;    16'd21123: out <= 16'h0312;
    16'd21124: out <= 16'hFFD4;    16'd21125: out <= 16'h01F1;    16'd21126: out <= 16'hFED4;    16'd21127: out <= 16'h0AC0;
    16'd21128: out <= 16'h0424;    16'd21129: out <= 16'h01CF;    16'd21130: out <= 16'h025B;    16'd21131: out <= 16'h0746;
    16'd21132: out <= 16'hFD93;    16'd21133: out <= 16'h03B1;    16'd21134: out <= 16'h03D0;    16'd21135: out <= 16'h0756;
    16'd21136: out <= 16'h0107;    16'd21137: out <= 16'hFFC1;    16'd21138: out <= 16'h0111;    16'd21139: out <= 16'hFEFB;
    16'd21140: out <= 16'h03AB;    16'd21141: out <= 16'h03C0;    16'd21142: out <= 16'h008D;    16'd21143: out <= 16'h057D;
    16'd21144: out <= 16'h0A83;    16'd21145: out <= 16'h00D0;    16'd21146: out <= 16'h0860;    16'd21147: out <= 16'h060D;
    16'd21148: out <= 16'h08F5;    16'd21149: out <= 16'h0226;    16'd21150: out <= 16'h080D;    16'd21151: out <= 16'h05A5;
    16'd21152: out <= 16'hFE58;    16'd21153: out <= 16'hFE19;    16'd21154: out <= 16'hFED9;    16'd21155: out <= 16'h0726;
    16'd21156: out <= 16'h0BDE;    16'd21157: out <= 16'hFC88;    16'd21158: out <= 16'hFF72;    16'd21159: out <= 16'h04BF;
    16'd21160: out <= 16'h03F0;    16'd21161: out <= 16'h0541;    16'd21162: out <= 16'h04E2;    16'd21163: out <= 16'h0745;
    16'd21164: out <= 16'h0216;    16'd21165: out <= 16'h042E;    16'd21166: out <= 16'h0B19;    16'd21167: out <= 16'h08F4;
    16'd21168: out <= 16'h06C2;    16'd21169: out <= 16'hFEC7;    16'd21170: out <= 16'h0659;    16'd21171: out <= 16'h0CCA;
    16'd21172: out <= 16'h0604;    16'd21173: out <= 16'h04BB;    16'd21174: out <= 16'h03F2;    16'd21175: out <= 16'hFFD3;
    16'd21176: out <= 16'h033C;    16'd21177: out <= 16'h06D3;    16'd21178: out <= 16'h06B6;    16'd21179: out <= 16'h018A;
    16'd21180: out <= 16'h032D;    16'd21181: out <= 16'h012C;    16'd21182: out <= 16'h0754;    16'd21183: out <= 16'h0B1B;
    16'd21184: out <= 16'h018D;    16'd21185: out <= 16'h0322;    16'd21186: out <= 16'h0820;    16'd21187: out <= 16'hFE1B;
    16'd21188: out <= 16'h0749;    16'd21189: out <= 16'hFBA8;    16'd21190: out <= 16'h07A5;    16'd21191: out <= 16'h048D;
    16'd21192: out <= 16'h016F;    16'd21193: out <= 16'h0326;    16'd21194: out <= 16'hFFAC;    16'd21195: out <= 16'hFE38;
    16'd21196: out <= 16'h0826;    16'd21197: out <= 16'h057E;    16'd21198: out <= 16'h0754;    16'd21199: out <= 16'h0236;
    16'd21200: out <= 16'h039E;    16'd21201: out <= 16'h02D5;    16'd21202: out <= 16'h05C6;    16'd21203: out <= 16'hFFE2;
    16'd21204: out <= 16'h00C6;    16'd21205: out <= 16'h04A1;    16'd21206: out <= 16'h07B8;    16'd21207: out <= 16'h0705;
    16'd21208: out <= 16'h030A;    16'd21209: out <= 16'h04AE;    16'd21210: out <= 16'hFC0E;    16'd21211: out <= 16'hFBEB;
    16'd21212: out <= 16'h0081;    16'd21213: out <= 16'hFEE4;    16'd21214: out <= 16'hFE2D;    16'd21215: out <= 16'h013F;
    16'd21216: out <= 16'h02F5;    16'd21217: out <= 16'h0363;    16'd21218: out <= 16'hF8FB;    16'd21219: out <= 16'h001B;
    16'd21220: out <= 16'h0273;    16'd21221: out <= 16'hFC2C;    16'd21222: out <= 16'h06CA;    16'd21223: out <= 16'h04CC;
    16'd21224: out <= 16'h029D;    16'd21225: out <= 16'hFD7F;    16'd21226: out <= 16'hFF2F;    16'd21227: out <= 16'h00F2;
    16'd21228: out <= 16'hF845;    16'd21229: out <= 16'h052B;    16'd21230: out <= 16'h0972;    16'd21231: out <= 16'hFF8B;
    16'd21232: out <= 16'hFF78;    16'd21233: out <= 16'hFCB7;    16'd21234: out <= 16'h01B6;    16'd21235: out <= 16'h01CB;
    16'd21236: out <= 16'h04EA;    16'd21237: out <= 16'hFCD3;    16'd21238: out <= 16'h070E;    16'd21239: out <= 16'hFFED;
    16'd21240: out <= 16'h022B;    16'd21241: out <= 16'hFED4;    16'd21242: out <= 16'hF9AC;    16'd21243: out <= 16'h0570;
    16'd21244: out <= 16'h03FA;    16'd21245: out <= 16'hFD76;    16'd21246: out <= 16'h001A;    16'd21247: out <= 16'h056A;
    16'd21248: out <= 16'h0554;    16'd21249: out <= 16'h0119;    16'd21250: out <= 16'h02AA;    16'd21251: out <= 16'hF9F1;
    16'd21252: out <= 16'hFB15;    16'd21253: out <= 16'hF7F4;    16'd21254: out <= 16'hFF3F;    16'd21255: out <= 16'h048B;
    16'd21256: out <= 16'h0239;    16'd21257: out <= 16'hF9FD;    16'd21258: out <= 16'hFC90;    16'd21259: out <= 16'hFA1C;
    16'd21260: out <= 16'hFB84;    16'd21261: out <= 16'h070E;    16'd21262: out <= 16'hFA46;    16'd21263: out <= 16'h04AA;
    16'd21264: out <= 16'h01EB;    16'd21265: out <= 16'hFF20;    16'd21266: out <= 16'h08D5;    16'd21267: out <= 16'h02BE;
    16'd21268: out <= 16'hFBD0;    16'd21269: out <= 16'h023D;    16'd21270: out <= 16'hFF8D;    16'd21271: out <= 16'hFB15;
    16'd21272: out <= 16'h0188;    16'd21273: out <= 16'h084D;    16'd21274: out <= 16'h0181;    16'd21275: out <= 16'h01FF;
    16'd21276: out <= 16'h0535;    16'd21277: out <= 16'h040B;    16'd21278: out <= 16'h0C86;    16'd21279: out <= 16'h0242;
    16'd21280: out <= 16'h0677;    16'd21281: out <= 16'hFAB9;    16'd21282: out <= 16'h01D5;    16'd21283: out <= 16'h0938;
    16'd21284: out <= 16'h0508;    16'd21285: out <= 16'h028B;    16'd21286: out <= 16'h04D4;    16'd21287: out <= 16'h03ED;
    16'd21288: out <= 16'h059C;    16'd21289: out <= 16'h0791;    16'd21290: out <= 16'h07B7;    16'd21291: out <= 16'h080F;
    16'd21292: out <= 16'h0275;    16'd21293: out <= 16'h0229;    16'd21294: out <= 16'h024F;    16'd21295: out <= 16'h01C3;
    16'd21296: out <= 16'h060F;    16'd21297: out <= 16'h04C6;    16'd21298: out <= 16'hFFDD;    16'd21299: out <= 16'h059F;
    16'd21300: out <= 16'hFC6C;    16'd21301: out <= 16'hFA51;    16'd21302: out <= 16'h03C3;    16'd21303: out <= 16'h033B;
    16'd21304: out <= 16'h0C44;    16'd21305: out <= 16'h0745;    16'd21306: out <= 16'h0066;    16'd21307: out <= 16'h04AF;
    16'd21308: out <= 16'h0014;    16'd21309: out <= 16'h096C;    16'd21310: out <= 16'h09BC;    16'd21311: out <= 16'h0096;
    16'd21312: out <= 16'h05A7;    16'd21313: out <= 16'hFD45;    16'd21314: out <= 16'hFF8F;    16'd21315: out <= 16'h0729;
    16'd21316: out <= 16'h064A;    16'd21317: out <= 16'h07F8;    16'd21318: out <= 16'hFF75;    16'd21319: out <= 16'h0522;
    16'd21320: out <= 16'h018E;    16'd21321: out <= 16'h0596;    16'd21322: out <= 16'h025D;    16'd21323: out <= 16'h05DC;
    16'd21324: out <= 16'hFCBB;    16'd21325: out <= 16'h0009;    16'd21326: out <= 16'h0180;    16'd21327: out <= 16'h03B0;
    16'd21328: out <= 16'hFB4C;    16'd21329: out <= 16'h0714;    16'd21330: out <= 16'hFDFE;    16'd21331: out <= 16'hFE93;
    16'd21332: out <= 16'h04C7;    16'd21333: out <= 16'h00BF;    16'd21334: out <= 16'h0295;    16'd21335: out <= 16'h0303;
    16'd21336: out <= 16'h0754;    16'd21337: out <= 16'h05EE;    16'd21338: out <= 16'h0BCE;    16'd21339: out <= 16'h01D8;
    16'd21340: out <= 16'h0750;    16'd21341: out <= 16'h04C9;    16'd21342: out <= 16'h0B7E;    16'd21343: out <= 16'h0118;
    16'd21344: out <= 16'h0182;    16'd21345: out <= 16'h032D;    16'd21346: out <= 16'h0188;    16'd21347: out <= 16'h01DE;
    16'd21348: out <= 16'h09AB;    16'd21349: out <= 16'h03C6;    16'd21350: out <= 16'hFD8B;    16'd21351: out <= 16'h0F8B;
    16'd21352: out <= 16'h019E;    16'd21353: out <= 16'h0758;    16'd21354: out <= 16'h064A;    16'd21355: out <= 16'h0627;
    16'd21356: out <= 16'hFF25;    16'd21357: out <= 16'h070F;    16'd21358: out <= 16'h071F;    16'd21359: out <= 16'h0498;
    16'd21360: out <= 16'hFEB4;    16'd21361: out <= 16'h052A;    16'd21362: out <= 16'hFFA7;    16'd21363: out <= 16'h0576;
    16'd21364: out <= 16'h03E9;    16'd21365: out <= 16'h0638;    16'd21366: out <= 16'h0969;    16'd21367: out <= 16'h0A0C;
    16'd21368: out <= 16'hFE20;    16'd21369: out <= 16'h0738;    16'd21370: out <= 16'h0618;    16'd21371: out <= 16'h081B;
    16'd21372: out <= 16'h0634;    16'd21373: out <= 16'h0518;    16'd21374: out <= 16'h07A2;    16'd21375: out <= 16'hFFD4;
    16'd21376: out <= 16'h0142;    16'd21377: out <= 16'h03FA;    16'd21378: out <= 16'h064B;    16'd21379: out <= 16'h0559;
    16'd21380: out <= 16'h025B;    16'd21381: out <= 16'h08DA;    16'd21382: out <= 16'hFAC3;    16'd21383: out <= 16'h014B;
    16'd21384: out <= 16'h00BA;    16'd21385: out <= 16'hFF10;    16'd21386: out <= 16'h0809;    16'd21387: out <= 16'h01F6;
    16'd21388: out <= 16'hFE2E;    16'd21389: out <= 16'h07D8;    16'd21390: out <= 16'h01DB;    16'd21391: out <= 16'h06B5;
    16'd21392: out <= 16'hFA8D;    16'd21393: out <= 16'h0398;    16'd21394: out <= 16'h00C6;    16'd21395: out <= 16'h021E;
    16'd21396: out <= 16'h0842;    16'd21397: out <= 16'h0C22;    16'd21398: out <= 16'h0024;    16'd21399: out <= 16'h0390;
    16'd21400: out <= 16'h07FA;    16'd21401: out <= 16'h05D1;    16'd21402: out <= 16'h0CD6;    16'd21403: out <= 16'h09C7;
    16'd21404: out <= 16'h0233;    16'd21405: out <= 16'hFE91;    16'd21406: out <= 16'h084F;    16'd21407: out <= 16'hFA11;
    16'd21408: out <= 16'hFFE8;    16'd21409: out <= 16'hFA80;    16'd21410: out <= 16'hFE94;    16'd21411: out <= 16'h00F9;
    16'd21412: out <= 16'h077C;    16'd21413: out <= 16'h08F1;    16'd21414: out <= 16'h05B9;    16'd21415: out <= 16'h06D4;
    16'd21416: out <= 16'hFEF4;    16'd21417: out <= 16'h0860;    16'd21418: out <= 16'h0172;    16'd21419: out <= 16'h0BDA;
    16'd21420: out <= 16'h04C8;    16'd21421: out <= 16'h080F;    16'd21422: out <= 16'hFEB8;    16'd21423: out <= 16'h03D1;
    16'd21424: out <= 16'h06E4;    16'd21425: out <= 16'h05B6;    16'd21426: out <= 16'h04BB;    16'd21427: out <= 16'h08F8;
    16'd21428: out <= 16'hFF15;    16'd21429: out <= 16'h0258;    16'd21430: out <= 16'h0263;    16'd21431: out <= 16'h086F;
    16'd21432: out <= 16'h0315;    16'd21433: out <= 16'h07C2;    16'd21434: out <= 16'h012D;    16'd21435: out <= 16'h0040;
    16'd21436: out <= 16'hFCCA;    16'd21437: out <= 16'h014D;    16'd21438: out <= 16'hFFA3;    16'd21439: out <= 16'h047C;
    16'd21440: out <= 16'h0751;    16'd21441: out <= 16'h035D;    16'd21442: out <= 16'h0518;    16'd21443: out <= 16'h04A7;
    16'd21444: out <= 16'h02FE;    16'd21445: out <= 16'h06CA;    16'd21446: out <= 16'h0468;    16'd21447: out <= 16'h0481;
    16'd21448: out <= 16'h04A2;    16'd21449: out <= 16'h068F;    16'd21450: out <= 16'h0342;    16'd21451: out <= 16'hFBE0;
    16'd21452: out <= 16'h039A;    16'd21453: out <= 16'h0759;    16'd21454: out <= 16'hFF6B;    16'd21455: out <= 16'hFFC7;
    16'd21456: out <= 16'h0736;    16'd21457: out <= 16'hFF98;    16'd21458: out <= 16'h06E9;    16'd21459: out <= 16'h07EA;
    16'd21460: out <= 16'h01E1;    16'd21461: out <= 16'h012E;    16'd21462: out <= 16'h0984;    16'd21463: out <= 16'h0347;
    16'd21464: out <= 16'h02E6;    16'd21465: out <= 16'hFF9A;    16'd21466: out <= 16'hFE84;    16'd21467: out <= 16'h0120;
    16'd21468: out <= 16'h0B00;    16'd21469: out <= 16'h051C;    16'd21470: out <= 16'h0169;    16'd21471: out <= 16'h03A1;
    16'd21472: out <= 16'h00D2;    16'd21473: out <= 16'hFB14;    16'd21474: out <= 16'hFC3B;    16'd21475: out <= 16'h0088;
    16'd21476: out <= 16'h0016;    16'd21477: out <= 16'h02D3;    16'd21478: out <= 16'hFC35;    16'd21479: out <= 16'hFE7B;
    16'd21480: out <= 16'h01F5;    16'd21481: out <= 16'h05A9;    16'd21482: out <= 16'h052D;    16'd21483: out <= 16'hFD30;
    16'd21484: out <= 16'hFF83;    16'd21485: out <= 16'hFB56;    16'd21486: out <= 16'hFF6C;    16'd21487: out <= 16'h035A;
    16'd21488: out <= 16'h05A1;    16'd21489: out <= 16'hFC03;    16'd21490: out <= 16'hFF7F;    16'd21491: out <= 16'hFDAB;
    16'd21492: out <= 16'h04FA;    16'd21493: out <= 16'h0129;    16'd21494: out <= 16'h006F;    16'd21495: out <= 16'hFDE5;
    16'd21496: out <= 16'h0630;    16'd21497: out <= 16'h0171;    16'd21498: out <= 16'hF78B;    16'd21499: out <= 16'hFCEA;
    16'd21500: out <= 16'h04A3;    16'd21501: out <= 16'hF7ED;    16'd21502: out <= 16'h079A;    16'd21503: out <= 16'h063E;
    16'd21504: out <= 16'h0955;    16'd21505: out <= 16'hFEFC;    16'd21506: out <= 16'hFDE7;    16'd21507: out <= 16'hF8B0;
    16'd21508: out <= 16'h03E4;    16'd21509: out <= 16'hFE27;    16'd21510: out <= 16'h0016;    16'd21511: out <= 16'h0084;
    16'd21512: out <= 16'hFD2D;    16'd21513: out <= 16'h04CB;    16'd21514: out <= 16'hFA2C;    16'd21515: out <= 16'h013D;
    16'd21516: out <= 16'h04C4;    16'd21517: out <= 16'h0345;    16'd21518: out <= 16'hFDBE;    16'd21519: out <= 16'h034B;
    16'd21520: out <= 16'hFAFC;    16'd21521: out <= 16'hFA6E;    16'd21522: out <= 16'hFCDA;    16'd21523: out <= 16'h0125;
    16'd21524: out <= 16'hFDAC;    16'd21525: out <= 16'hFFA2;    16'd21526: out <= 16'h0067;    16'd21527: out <= 16'hFDB3;
    16'd21528: out <= 16'h00E2;    16'd21529: out <= 16'h02DE;    16'd21530: out <= 16'hFE36;    16'd21531: out <= 16'h00F9;
    16'd21532: out <= 16'h08B5;    16'd21533: out <= 16'h0A8B;    16'd21534: out <= 16'h022D;    16'd21535: out <= 16'hFAAC;
    16'd21536: out <= 16'h0553;    16'd21537: out <= 16'h0239;    16'd21538: out <= 16'h022E;    16'd21539: out <= 16'h065B;
    16'd21540: out <= 16'hFF68;    16'd21541: out <= 16'h003B;    16'd21542: out <= 16'h0777;    16'd21543: out <= 16'h069B;
    16'd21544: out <= 16'h080E;    16'd21545: out <= 16'h09D0;    16'd21546: out <= 16'h0579;    16'd21547: out <= 16'h01D5;
    16'd21548: out <= 16'h072D;    16'd21549: out <= 16'h07D9;    16'd21550: out <= 16'h0082;    16'd21551: out <= 16'hFE99;
    16'd21552: out <= 16'h07A6;    16'd21553: out <= 16'h0976;    16'd21554: out <= 16'h0065;    16'd21555: out <= 16'h0500;
    16'd21556: out <= 16'hFEB3;    16'd21557: out <= 16'h0142;    16'd21558: out <= 16'h0313;    16'd21559: out <= 16'h03A6;
    16'd21560: out <= 16'hFEA6;    16'd21561: out <= 16'hFEBF;    16'd21562: out <= 16'h05C5;    16'd21563: out <= 16'hF938;
    16'd21564: out <= 16'h04FF;    16'd21565: out <= 16'h0A7A;    16'd21566: out <= 16'h0000;    16'd21567: out <= 16'h026D;
    16'd21568: out <= 16'hFC4E;    16'd21569: out <= 16'h0641;    16'd21570: out <= 16'h0179;    16'd21571: out <= 16'h013F;
    16'd21572: out <= 16'h0B41;    16'd21573: out <= 16'hFEEC;    16'd21574: out <= 16'hFEA3;    16'd21575: out <= 16'h0A73;
    16'd21576: out <= 16'h075E;    16'd21577: out <= 16'h0217;    16'd21578: out <= 16'h03DC;    16'd21579: out <= 16'h05DD;
    16'd21580: out <= 16'h079E;    16'd21581: out <= 16'h03C5;    16'd21582: out <= 16'hFCB5;    16'd21583: out <= 16'h0102;
    16'd21584: out <= 16'h0237;    16'd21585: out <= 16'hFD77;    16'd21586: out <= 16'hFC89;    16'd21587: out <= 16'hFDE4;
    16'd21588: out <= 16'h0263;    16'd21589: out <= 16'hFDA8;    16'd21590: out <= 16'h0630;    16'd21591: out <= 16'h0545;
    16'd21592: out <= 16'h059C;    16'd21593: out <= 16'h07FA;    16'd21594: out <= 16'h0274;    16'd21595: out <= 16'h0830;
    16'd21596: out <= 16'h003D;    16'd21597: out <= 16'h0160;    16'd21598: out <= 16'h0087;    16'd21599: out <= 16'h0417;
    16'd21600: out <= 16'h0701;    16'd21601: out <= 16'h06AB;    16'd21602: out <= 16'hFC9A;    16'd21603: out <= 16'hFCC4;
    16'd21604: out <= 16'h068C;    16'd21605: out <= 16'h007B;    16'd21606: out <= 16'h03FC;    16'd21607: out <= 16'h0727;
    16'd21608: out <= 16'h0654;    16'd21609: out <= 16'h04D0;    16'd21610: out <= 16'h019B;    16'd21611: out <= 16'h08F8;
    16'd21612: out <= 16'h0757;    16'd21613: out <= 16'h04B7;    16'd21614: out <= 16'h0264;    16'd21615: out <= 16'h01BA;
    16'd21616: out <= 16'h05B9;    16'd21617: out <= 16'h05FA;    16'd21618: out <= 16'hFFD1;    16'd21619: out <= 16'h011E;
    16'd21620: out <= 16'h0872;    16'd21621: out <= 16'h01C4;    16'd21622: out <= 16'h069D;    16'd21623: out <= 16'h0931;
    16'd21624: out <= 16'h0469;    16'd21625: out <= 16'h07EF;    16'd21626: out <= 16'h0050;    16'd21627: out <= 16'h04D8;
    16'd21628: out <= 16'h0134;    16'd21629: out <= 16'h04F9;    16'd21630: out <= 16'h0C10;    16'd21631: out <= 16'h0436;
    16'd21632: out <= 16'h05BE;    16'd21633: out <= 16'h05F1;    16'd21634: out <= 16'h04F1;    16'd21635: out <= 16'h0769;
    16'd21636: out <= 16'h031E;    16'd21637: out <= 16'h0710;    16'd21638: out <= 16'h04A5;    16'd21639: out <= 16'h05FB;
    16'd21640: out <= 16'h0499;    16'd21641: out <= 16'h060B;    16'd21642: out <= 16'h068F;    16'd21643: out <= 16'h044F;
    16'd21644: out <= 16'h0AE7;    16'd21645: out <= 16'h0BF8;    16'd21646: out <= 16'h00F1;    16'd21647: out <= 16'h0702;
    16'd21648: out <= 16'hFF3B;    16'd21649: out <= 16'h06B2;    16'd21650: out <= 16'h0575;    16'd21651: out <= 16'hFF2A;
    16'd21652: out <= 16'h0813;    16'd21653: out <= 16'h0674;    16'd21654: out <= 16'h030D;    16'd21655: out <= 16'hFE58;
    16'd21656: out <= 16'h0173;    16'd21657: out <= 16'hFBD3;    16'd21658: out <= 16'hFE37;    16'd21659: out <= 16'hF67D;
    16'd21660: out <= 16'h0199;    16'd21661: out <= 16'h008B;    16'd21662: out <= 16'h0767;    16'd21663: out <= 16'h0236;
    16'd21664: out <= 16'hF82A;    16'd21665: out <= 16'hFBBC;    16'd21666: out <= 16'h0277;    16'd21667: out <= 16'hFF8A;
    16'd21668: out <= 16'h03A0;    16'd21669: out <= 16'hFCEF;    16'd21670: out <= 16'hFCDA;    16'd21671: out <= 16'hFDF7;
    16'd21672: out <= 16'h0A6F;    16'd21673: out <= 16'hF941;    16'd21674: out <= 16'h08B1;    16'd21675: out <= 16'hFB66;
    16'd21676: out <= 16'h0B57;    16'd21677: out <= 16'h0192;    16'd21678: out <= 16'h05B9;    16'd21679: out <= 16'h05FC;
    16'd21680: out <= 16'h006E;    16'd21681: out <= 16'h07C5;    16'd21682: out <= 16'h06CE;    16'd21683: out <= 16'h008C;
    16'd21684: out <= 16'h066D;    16'd21685: out <= 16'h0349;    16'd21686: out <= 16'h0212;    16'd21687: out <= 16'hFF60;
    16'd21688: out <= 16'h045D;    16'd21689: out <= 16'h0D25;    16'd21690: out <= 16'h0797;    16'd21691: out <= 16'h06A6;
    16'd21692: out <= 16'h0B01;    16'd21693: out <= 16'h043C;    16'd21694: out <= 16'h0460;    16'd21695: out <= 16'h0AC0;
    16'd21696: out <= 16'h04DD;    16'd21697: out <= 16'h0597;    16'd21698: out <= 16'h0787;    16'd21699: out <= 16'h0699;
    16'd21700: out <= 16'h0437;    16'd21701: out <= 16'hFD76;    16'd21702: out <= 16'h02C2;    16'd21703: out <= 16'h00BA;
    16'd21704: out <= 16'h0695;    16'd21705: out <= 16'h001B;    16'd21706: out <= 16'h04D0;    16'd21707: out <= 16'h01C6;
    16'd21708: out <= 16'hFF87;    16'd21709: out <= 16'h022A;    16'd21710: out <= 16'h0588;    16'd21711: out <= 16'hFFA9;
    16'd21712: out <= 16'h0848;    16'd21713: out <= 16'hFEF7;    16'd21714: out <= 16'h0452;    16'd21715: out <= 16'h04EB;
    16'd21716: out <= 16'h0214;    16'd21717: out <= 16'h0499;    16'd21718: out <= 16'h034A;    16'd21719: out <= 16'h0720;
    16'd21720: out <= 16'h01F7;    16'd21721: out <= 16'h0700;    16'd21722: out <= 16'hFFE4;    16'd21723: out <= 16'h0085;
    16'd21724: out <= 16'hFB9E;    16'd21725: out <= 16'h00E6;    16'd21726: out <= 16'hFE99;    16'd21727: out <= 16'h0180;
    16'd21728: out <= 16'hFD16;    16'd21729: out <= 16'h084F;    16'd21730: out <= 16'hFB9A;    16'd21731: out <= 16'h03E9;
    16'd21732: out <= 16'hFEB2;    16'd21733: out <= 16'hFD10;    16'd21734: out <= 16'h0205;    16'd21735: out <= 16'h0179;
    16'd21736: out <= 16'hFE5F;    16'd21737: out <= 16'h0358;    16'd21738: out <= 16'h0066;    16'd21739: out <= 16'h001A;
    16'd21740: out <= 16'hF895;    16'd21741: out <= 16'h077B;    16'd21742: out <= 16'hFF23;    16'd21743: out <= 16'h057E;
    16'd21744: out <= 16'h02C2;    16'd21745: out <= 16'hFBB1;    16'd21746: out <= 16'hFBB2;    16'd21747: out <= 16'hFF27;
    16'd21748: out <= 16'h082C;    16'd21749: out <= 16'hFE29;    16'd21750: out <= 16'h00BD;    16'd21751: out <= 16'h0123;
    16'd21752: out <= 16'hFDD9;    16'd21753: out <= 16'hFE12;    16'd21754: out <= 16'hFFEB;    16'd21755: out <= 16'h05B4;
    16'd21756: out <= 16'hFB72;    16'd21757: out <= 16'h005F;    16'd21758: out <= 16'hFF53;    16'd21759: out <= 16'hF97E;
    16'd21760: out <= 16'hFFBF;    16'd21761: out <= 16'hFDB7;    16'd21762: out <= 16'hFF9F;    16'd21763: out <= 16'hFF15;
    16'd21764: out <= 16'hFA4A;    16'd21765: out <= 16'h00F7;    16'd21766: out <= 16'h00E8;    16'd21767: out <= 16'h02F5;
    16'd21768: out <= 16'hFD56;    16'd21769: out <= 16'hFD94;    16'd21770: out <= 16'h0170;    16'd21771: out <= 16'h0607;
    16'd21772: out <= 16'hFCE5;    16'd21773: out <= 16'h0591;    16'd21774: out <= 16'hFF15;    16'd21775: out <= 16'hFE2F;
    16'd21776: out <= 16'h0430;    16'd21777: out <= 16'hFD19;    16'd21778: out <= 16'h073F;    16'd21779: out <= 16'hF3BE;
    16'd21780: out <= 16'h03D0;    16'd21781: out <= 16'h0095;    16'd21782: out <= 16'hFCF2;    16'd21783: out <= 16'h0149;
    16'd21784: out <= 16'h00EA;    16'd21785: out <= 16'h0664;    16'd21786: out <= 16'h0541;    16'd21787: out <= 16'hFD61;
    16'd21788: out <= 16'h0A15;    16'd21789: out <= 16'h04EB;    16'd21790: out <= 16'h06B6;    16'd21791: out <= 16'h07F1;
    16'd21792: out <= 16'h05DA;    16'd21793: out <= 16'h049D;    16'd21794: out <= 16'h0341;    16'd21795: out <= 16'h0783;
    16'd21796: out <= 16'hF942;    16'd21797: out <= 16'h06E3;    16'd21798: out <= 16'h0447;    16'd21799: out <= 16'h05C9;
    16'd21800: out <= 16'h04E0;    16'd21801: out <= 16'h05A0;    16'd21802: out <= 16'h03D7;    16'd21803: out <= 16'h051B;
    16'd21804: out <= 16'h0C6A;    16'd21805: out <= 16'h0CEC;    16'd21806: out <= 16'h060E;    16'd21807: out <= 16'h029C;
    16'd21808: out <= 16'h0355;    16'd21809: out <= 16'h0825;    16'd21810: out <= 16'h0419;    16'd21811: out <= 16'h0467;
    16'd21812: out <= 16'h012E;    16'd21813: out <= 16'hFECE;    16'd21814: out <= 16'hFE78;    16'd21815: out <= 16'h0074;
    16'd21816: out <= 16'h07A0;    16'd21817: out <= 16'h01BA;    16'd21818: out <= 16'h045D;    16'd21819: out <= 16'h000E;
    16'd21820: out <= 16'h059D;    16'd21821: out <= 16'h061A;    16'd21822: out <= 16'h051C;    16'd21823: out <= 16'h01B2;
    16'd21824: out <= 16'h0607;    16'd21825: out <= 16'h0334;    16'd21826: out <= 16'h093F;    16'd21827: out <= 16'hFD06;
    16'd21828: out <= 16'h044A;    16'd21829: out <= 16'hFF6D;    16'd21830: out <= 16'h0450;    16'd21831: out <= 16'h0918;
    16'd21832: out <= 16'h05D5;    16'd21833: out <= 16'h042A;    16'd21834: out <= 16'h06E0;    16'd21835: out <= 16'h022F;
    16'd21836: out <= 16'h071A;    16'd21837: out <= 16'hFD24;    16'd21838: out <= 16'h03DA;    16'd21839: out <= 16'hFFB9;
    16'd21840: out <= 16'hFD4D;    16'd21841: out <= 16'h04C4;    16'd21842: out <= 16'h0354;    16'd21843: out <= 16'h02F5;
    16'd21844: out <= 16'h0214;    16'd21845: out <= 16'h091A;    16'd21846: out <= 16'h032A;    16'd21847: out <= 16'h068F;
    16'd21848: out <= 16'h0529;    16'd21849: out <= 16'h0569;    16'd21850: out <= 16'h08A4;    16'd21851: out <= 16'h0453;
    16'd21852: out <= 16'h07AC;    16'd21853: out <= 16'h0608;    16'd21854: out <= 16'h0419;    16'd21855: out <= 16'h097F;
    16'd21856: out <= 16'h041E;    16'd21857: out <= 16'h06C2;    16'd21858: out <= 16'h0919;    16'd21859: out <= 16'h053D;
    16'd21860: out <= 16'h0269;    16'd21861: out <= 16'h07D1;    16'd21862: out <= 16'h05CF;    16'd21863: out <= 16'h09C0;
    16'd21864: out <= 16'hFD89;    16'd21865: out <= 16'h074B;    16'd21866: out <= 16'h047F;    16'd21867: out <= 16'hFAAB;
    16'd21868: out <= 16'h0B7F;    16'd21869: out <= 16'h00A6;    16'd21870: out <= 16'h0713;    16'd21871: out <= 16'h0727;
    16'd21872: out <= 16'h07F7;    16'd21873: out <= 16'h0102;    16'd21874: out <= 16'h01C2;    16'd21875: out <= 16'h048D;
    16'd21876: out <= 16'h0264;    16'd21877: out <= 16'h03C7;    16'd21878: out <= 16'hFEFB;    16'd21879: out <= 16'hFF6C;
    16'd21880: out <= 16'h0239;    16'd21881: out <= 16'h017D;    16'd21882: out <= 16'h0255;    16'd21883: out <= 16'h0253;
    16'd21884: out <= 16'h02FE;    16'd21885: out <= 16'h02D0;    16'd21886: out <= 16'h0ABB;    16'd21887: out <= 16'h0427;
    16'd21888: out <= 16'h0420;    16'd21889: out <= 16'h0BC0;    16'd21890: out <= 16'h01E2;    16'd21891: out <= 16'hFB3D;
    16'd21892: out <= 16'hFEC9;    16'd21893: out <= 16'h073F;    16'd21894: out <= 16'h0445;    16'd21895: out <= 16'h00B2;
    16'd21896: out <= 16'h06EB;    16'd21897: out <= 16'h056F;    16'd21898: out <= 16'hFED1;    16'd21899: out <= 16'h0190;
    16'd21900: out <= 16'h0172;    16'd21901: out <= 16'h04A2;    16'd21902: out <= 16'h0B1F;    16'd21903: out <= 16'h0323;
    16'd21904: out <= 16'hFED3;    16'd21905: out <= 16'h0697;    16'd21906: out <= 16'hFFB1;    16'd21907: out <= 16'h0413;
    16'd21908: out <= 16'h0292;    16'd21909: out <= 16'h035F;    16'd21910: out <= 16'h07EE;    16'd21911: out <= 16'h09B1;
    16'd21912: out <= 16'h0196;    16'd21913: out <= 16'h0005;    16'd21914: out <= 16'hFE47;    16'd21915: out <= 16'hFCD9;
    16'd21916: out <= 16'hFC67;    16'd21917: out <= 16'hFDFE;    16'd21918: out <= 16'hFF3C;    16'd21919: out <= 16'hFE7A;
    16'd21920: out <= 16'hFC7E;    16'd21921: out <= 16'h0421;    16'd21922: out <= 16'h0471;    16'd21923: out <= 16'h0144;
    16'd21924: out <= 16'h0054;    16'd21925: out <= 16'h0480;    16'd21926: out <= 16'h00C7;    16'd21927: out <= 16'h0504;
    16'd21928: out <= 16'h07BB;    16'd21929: out <= 16'h037C;    16'd21930: out <= 16'h03B5;    16'd21931: out <= 16'h0485;
    16'd21932: out <= 16'hFB3E;    16'd21933: out <= 16'h04EE;    16'd21934: out <= 16'h02C8;    16'd21935: out <= 16'h083B;
    16'd21936: out <= 16'hFF30;    16'd21937: out <= 16'h0300;    16'd21938: out <= 16'h029B;    16'd21939: out <= 16'h0ABC;
    16'd21940: out <= 16'h0433;    16'd21941: out <= 16'h0977;    16'd21942: out <= 16'h07A6;    16'd21943: out <= 16'h035B;
    16'd21944: out <= 16'h0436;    16'd21945: out <= 16'h04E9;    16'd21946: out <= 16'h0714;    16'd21947: out <= 16'hFF68;
    16'd21948: out <= 16'h02A5;    16'd21949: out <= 16'h0215;    16'd21950: out <= 16'h0361;    16'd21951: out <= 16'h04F3;
    16'd21952: out <= 16'hFC9C;    16'd21953: out <= 16'hFEC2;    16'd21954: out <= 16'hFC54;    16'd21955: out <= 16'hFDAE;
    16'd21956: out <= 16'h06D1;    16'd21957: out <= 16'hFC2B;    16'd21958: out <= 16'h0A25;    16'd21959: out <= 16'hFAE9;
    16'd21960: out <= 16'h052C;    16'd21961: out <= 16'h0434;    16'd21962: out <= 16'h03E1;    16'd21963: out <= 16'h056B;
    16'd21964: out <= 16'h0197;    16'd21965: out <= 16'h0092;    16'd21966: out <= 16'hFC6E;    16'd21967: out <= 16'h0400;
    16'd21968: out <= 16'h0217;    16'd21969: out <= 16'h0134;    16'd21970: out <= 16'h0189;    16'd21971: out <= 16'h00C3;
    16'd21972: out <= 16'h06ED;    16'd21973: out <= 16'h027E;    16'd21974: out <= 16'h0D19;    16'd21975: out <= 16'hFE29;
    16'd21976: out <= 16'h02A8;    16'd21977: out <= 16'h01ED;    16'd21978: out <= 16'hFD22;    16'd21979: out <= 16'hFBF1;
    16'd21980: out <= 16'h024A;    16'd21981: out <= 16'h0033;    16'd21982: out <= 16'hFEE9;    16'd21983: out <= 16'h0123;
    16'd21984: out <= 16'h00A0;    16'd21985: out <= 16'hFCE7;    16'd21986: out <= 16'h051C;    16'd21987: out <= 16'h0043;
    16'd21988: out <= 16'hFF5A;    16'd21989: out <= 16'h02DF;    16'd21990: out <= 16'h01BA;    16'd21991: out <= 16'h03A1;
    16'd21992: out <= 16'hFD11;    16'd21993: out <= 16'hFF80;    16'd21994: out <= 16'h02F4;    16'd21995: out <= 16'h03BE;
    16'd21996: out <= 16'h0113;    16'd21997: out <= 16'h0205;    16'd21998: out <= 16'hFDC8;    16'd21999: out <= 16'hFA25;
    16'd22000: out <= 16'h0583;    16'd22001: out <= 16'hFB16;    16'd22002: out <= 16'hFF61;    16'd22003: out <= 16'h04ED;
    16'd22004: out <= 16'h01A7;    16'd22005: out <= 16'hFF4D;    16'd22006: out <= 16'h0A5F;    16'd22007: out <= 16'hFCEF;
    16'd22008: out <= 16'hFB2A;    16'd22009: out <= 16'h0268;    16'd22010: out <= 16'hFD91;    16'd22011: out <= 16'hFC2B;
    16'd22012: out <= 16'h0171;    16'd22013: out <= 16'h020D;    16'd22014: out <= 16'h013C;    16'd22015: out <= 16'hFDCA;
    16'd22016: out <= 16'hFEF8;    16'd22017: out <= 16'h027E;    16'd22018: out <= 16'h0241;    16'd22019: out <= 16'h0434;
    16'd22020: out <= 16'h0445;    16'd22021: out <= 16'hFAA8;    16'd22022: out <= 16'h01A1;    16'd22023: out <= 16'hFE6C;
    16'd22024: out <= 16'h0533;    16'd22025: out <= 16'h0640;    16'd22026: out <= 16'hFCC0;    16'd22027: out <= 16'h030D;
    16'd22028: out <= 16'h0385;    16'd22029: out <= 16'hF97C;    16'd22030: out <= 16'hFFBE;    16'd22031: out <= 16'hFAAF;
    16'd22032: out <= 16'h0380;    16'd22033: out <= 16'h01AB;    16'd22034: out <= 16'hFF67;    16'd22035: out <= 16'h0491;
    16'd22036: out <= 16'hF8F2;    16'd22037: out <= 16'h0037;    16'd22038: out <= 16'h045B;    16'd22039: out <= 16'h0105;
    16'd22040: out <= 16'hFBC4;    16'd22041: out <= 16'h066A;    16'd22042: out <= 16'h0392;    16'd22043: out <= 16'h014B;
    16'd22044: out <= 16'h0047;    16'd22045: out <= 16'h0057;    16'd22046: out <= 16'h05BC;    16'd22047: out <= 16'h01E5;
    16'd22048: out <= 16'h0662;    16'd22049: out <= 16'h06E4;    16'd22050: out <= 16'h07F2;    16'd22051: out <= 16'hFDF9;
    16'd22052: out <= 16'hFDD1;    16'd22053: out <= 16'h02AB;    16'd22054: out <= 16'h075A;    16'd22055: out <= 16'h0706;
    16'd22056: out <= 16'h0072;    16'd22057: out <= 16'h049F;    16'd22058: out <= 16'h0351;    16'd22059: out <= 16'h02F1;
    16'd22060: out <= 16'h0269;    16'd22061: out <= 16'h002B;    16'd22062: out <= 16'h0878;    16'd22063: out <= 16'h0644;
    16'd22064: out <= 16'hFD0E;    16'd22065: out <= 16'h0D10;    16'd22066: out <= 16'h1197;    16'd22067: out <= 16'h06BF;
    16'd22068: out <= 16'h0ABF;    16'd22069: out <= 16'h01DB;    16'd22070: out <= 16'h043C;    16'd22071: out <= 16'h063D;
    16'd22072: out <= 16'h09E6;    16'd22073: out <= 16'h0442;    16'd22074: out <= 16'h0984;    16'd22075: out <= 16'hFFA6;
    16'd22076: out <= 16'h094B;    16'd22077: out <= 16'hF98E;    16'd22078: out <= 16'h063D;    16'd22079: out <= 16'h03E2;
    16'd22080: out <= 16'h0760;    16'd22081: out <= 16'h04ED;    16'd22082: out <= 16'h02A3;    16'd22083: out <= 16'h07E1;
    16'd22084: out <= 16'hFCD2;    16'd22085: out <= 16'hFF79;    16'd22086: out <= 16'hFF4F;    16'd22087: out <= 16'h076E;
    16'd22088: out <= 16'h0740;    16'd22089: out <= 16'h0758;    16'd22090: out <= 16'h0857;    16'd22091: out <= 16'h07AB;
    16'd22092: out <= 16'hFFD7;    16'd22093: out <= 16'hFC20;    16'd22094: out <= 16'h0783;    16'd22095: out <= 16'h01DB;
    16'd22096: out <= 16'hFD57;    16'd22097: out <= 16'h0620;    16'd22098: out <= 16'hFFBF;    16'd22099: out <= 16'h023B;
    16'd22100: out <= 16'h0356;    16'd22101: out <= 16'h01CD;    16'd22102: out <= 16'h0608;    16'd22103: out <= 16'h0B0E;
    16'd22104: out <= 16'h0519;    16'd22105: out <= 16'h05E4;    16'd22106: out <= 16'h0CCD;    16'd22107: out <= 16'h0097;
    16'd22108: out <= 16'h0107;    16'd22109: out <= 16'h08DF;    16'd22110: out <= 16'hFF20;    16'd22111: out <= 16'hFF5F;
    16'd22112: out <= 16'hFFF9;    16'd22113: out <= 16'h077B;    16'd22114: out <= 16'h0235;    16'd22115: out <= 16'h0620;
    16'd22116: out <= 16'h0158;    16'd22117: out <= 16'h005C;    16'd22118: out <= 16'hFEB5;    16'd22119: out <= 16'h06F7;
    16'd22120: out <= 16'h03DE;    16'd22121: out <= 16'h0745;    16'd22122: out <= 16'hFD0B;    16'd22123: out <= 16'h0309;
    16'd22124: out <= 16'h0BC8;    16'd22125: out <= 16'h022C;    16'd22126: out <= 16'h00D8;    16'd22127: out <= 16'h0196;
    16'd22128: out <= 16'h05E2;    16'd22129: out <= 16'h0609;    16'd22130: out <= 16'h0563;    16'd22131: out <= 16'h02E7;
    16'd22132: out <= 16'h0540;    16'd22133: out <= 16'h0211;    16'd22134: out <= 16'h0310;    16'd22135: out <= 16'h09E9;
    16'd22136: out <= 16'h02A1;    16'd22137: out <= 16'h044C;    16'd22138: out <= 16'hFF33;    16'd22139: out <= 16'hFD39;
    16'd22140: out <= 16'h0023;    16'd22141: out <= 16'hFF68;    16'd22142: out <= 16'h0782;    16'd22143: out <= 16'h0436;
    16'd22144: out <= 16'h099B;    16'd22145: out <= 16'hFBFD;    16'd22146: out <= 16'h0792;    16'd22147: out <= 16'h04EF;
    16'd22148: out <= 16'h0911;    16'd22149: out <= 16'h03BD;    16'd22150: out <= 16'h077E;    16'd22151: out <= 16'hFED9;
    16'd22152: out <= 16'h0274;    16'd22153: out <= 16'h013C;    16'd22154: out <= 16'h0745;    16'd22155: out <= 16'hFD7D;
    16'd22156: out <= 16'h0008;    16'd22157: out <= 16'h03EF;    16'd22158: out <= 16'h0848;    16'd22159: out <= 16'h07B6;
    16'd22160: out <= 16'h003F;    16'd22161: out <= 16'h0119;    16'd22162: out <= 16'h0148;    16'd22163: out <= 16'h0480;
    16'd22164: out <= 16'h05FA;    16'd22165: out <= 16'h00F5;    16'd22166: out <= 16'h00D1;    16'd22167: out <= 16'hFB91;
    16'd22168: out <= 16'hFE84;    16'd22169: out <= 16'h003A;    16'd22170: out <= 16'h03D5;    16'd22171: out <= 16'h0549;
    16'd22172: out <= 16'hFF0F;    16'd22173: out <= 16'h0208;    16'd22174: out <= 16'hFAED;    16'd22175: out <= 16'hFC00;
    16'd22176: out <= 16'hFF88;    16'd22177: out <= 16'h02E6;    16'd22178: out <= 16'h05B8;    16'd22179: out <= 16'hF9BA;
    16'd22180: out <= 16'hFE64;    16'd22181: out <= 16'hFD99;    16'd22182: out <= 16'h08AA;    16'd22183: out <= 16'h0387;
    16'd22184: out <= 16'h024F;    16'd22185: out <= 16'h04B6;    16'd22186: out <= 16'h01BC;    16'd22187: out <= 16'h01DB;
    16'd22188: out <= 16'h0A2B;    16'd22189: out <= 16'h07F4;    16'd22190: out <= 16'h03B4;    16'd22191: out <= 16'h0597;
    16'd22192: out <= 16'h0576;    16'd22193: out <= 16'h0A2D;    16'd22194: out <= 16'h09B9;    16'd22195: out <= 16'h0CDA;
    16'd22196: out <= 16'h05D2;    16'd22197: out <= 16'h0715;    16'd22198: out <= 16'h01F3;    16'd22199: out <= 16'h03CF;
    16'd22200: out <= 16'h0BA8;    16'd22201: out <= 16'h0406;    16'd22202: out <= 16'h08AF;    16'd22203: out <= 16'h06B9;
    16'd22204: out <= 16'h00D4;    16'd22205: out <= 16'h054B;    16'd22206: out <= 16'h05FC;    16'd22207: out <= 16'h08FA;
    16'd22208: out <= 16'h0019;    16'd22209: out <= 16'hFE17;    16'd22210: out <= 16'h0929;    16'd22211: out <= 16'h0786;
    16'd22212: out <= 16'h0377;    16'd22213: out <= 16'h027E;    16'd22214: out <= 16'h0182;    16'd22215: out <= 16'hFF03;
    16'd22216: out <= 16'h0485;    16'd22217: out <= 16'h0416;    16'd22218: out <= 16'h04F5;    16'd22219: out <= 16'h027C;
    16'd22220: out <= 16'hFCB0;    16'd22221: out <= 16'h0239;    16'd22222: out <= 16'h008A;    16'd22223: out <= 16'h053F;
    16'd22224: out <= 16'h0695;    16'd22225: out <= 16'h04E2;    16'd22226: out <= 16'h0160;    16'd22227: out <= 16'h019A;
    16'd22228: out <= 16'h0767;    16'd22229: out <= 16'hFE78;    16'd22230: out <= 16'h05F6;    16'd22231: out <= 16'h00D7;
    16'd22232: out <= 16'h04FD;    16'd22233: out <= 16'h0657;    16'd22234: out <= 16'hFE8B;    16'd22235: out <= 16'h0254;
    16'd22236: out <= 16'h0435;    16'd22237: out <= 16'h0148;    16'd22238: out <= 16'h0403;    16'd22239: out <= 16'h050F;
    16'd22240: out <= 16'hFE58;    16'd22241: out <= 16'h0594;    16'd22242: out <= 16'hFED6;    16'd22243: out <= 16'hFF09;
    16'd22244: out <= 16'h04BB;    16'd22245: out <= 16'h04D1;    16'd22246: out <= 16'hFF25;    16'd22247: out <= 16'hFA5D;
    16'd22248: out <= 16'hFE31;    16'd22249: out <= 16'hFD65;    16'd22250: out <= 16'h01B1;    16'd22251: out <= 16'h0364;
    16'd22252: out <= 16'hF8A8;    16'd22253: out <= 16'h0286;    16'd22254: out <= 16'h0451;    16'd22255: out <= 16'hFE0A;
    16'd22256: out <= 16'hFDAD;    16'd22257: out <= 16'hF88C;    16'd22258: out <= 16'h04FD;    16'd22259: out <= 16'h04CA;
    16'd22260: out <= 16'hFAF5;    16'd22261: out <= 16'hFE87;    16'd22262: out <= 16'hFF06;    16'd22263: out <= 16'h03F9;
    16'd22264: out <= 16'hF85D;    16'd22265: out <= 16'hFDC9;    16'd22266: out <= 16'h0242;    16'd22267: out <= 16'h03D1;
    16'd22268: out <= 16'h045A;    16'd22269: out <= 16'h051E;    16'd22270: out <= 16'h02BD;    16'd22271: out <= 16'h02AE;
    16'd22272: out <= 16'h0315;    16'd22273: out <= 16'hFD88;    16'd22274: out <= 16'hFD67;    16'd22275: out <= 16'hFF76;
    16'd22276: out <= 16'hFD7A;    16'd22277: out <= 16'h04DC;    16'd22278: out <= 16'h02FD;    16'd22279: out <= 16'hFDAA;
    16'd22280: out <= 16'hFF0A;    16'd22281: out <= 16'hFA6D;    16'd22282: out <= 16'hF6DF;    16'd22283: out <= 16'hFD35;
    16'd22284: out <= 16'h0AC2;    16'd22285: out <= 16'hFFFB;    16'd22286: out <= 16'hFD39;    16'd22287: out <= 16'hFD66;
    16'd22288: out <= 16'h015A;    16'd22289: out <= 16'h06C9;    16'd22290: out <= 16'h0282;    16'd22291: out <= 16'hFA1C;
    16'd22292: out <= 16'hF966;    16'd22293: out <= 16'hFD1F;    16'd22294: out <= 16'h0181;    16'd22295: out <= 16'h0302;
    16'd22296: out <= 16'hFD20;    16'd22297: out <= 16'h00DF;    16'd22298: out <= 16'h0519;    16'd22299: out <= 16'h026A;
    16'd22300: out <= 16'hFE7A;    16'd22301: out <= 16'h0406;    16'd22302: out <= 16'h06C0;    16'd22303: out <= 16'h071C;
    16'd22304: out <= 16'h051A;    16'd22305: out <= 16'h0A87;    16'd22306: out <= 16'h0409;    16'd22307: out <= 16'h0567;
    16'd22308: out <= 16'h03DC;    16'd22309: out <= 16'h03D6;    16'd22310: out <= 16'hFF4B;    16'd22311: out <= 16'hFE1B;
    16'd22312: out <= 16'h0B67;    16'd22313: out <= 16'h0258;    16'd22314: out <= 16'h02DF;    16'd22315: out <= 16'hFF1E;
    16'd22316: out <= 16'h0337;    16'd22317: out <= 16'h0DB8;    16'd22318: out <= 16'hFCD5;    16'd22319: out <= 16'hF9EE;
    16'd22320: out <= 16'h00BB;    16'd22321: out <= 16'h0209;    16'd22322: out <= 16'h063B;    16'd22323: out <= 16'h09B9;
    16'd22324: out <= 16'h0506;    16'd22325: out <= 16'h0488;    16'd22326: out <= 16'h0723;    16'd22327: out <= 16'hFF04;
    16'd22328: out <= 16'hFDCD;    16'd22329: out <= 16'hFD0E;    16'd22330: out <= 16'h079E;    16'd22331: out <= 16'h08C6;
    16'd22332: out <= 16'h0A72;    16'd22333: out <= 16'h071D;    16'd22334: out <= 16'h00F9;    16'd22335: out <= 16'h055B;
    16'd22336: out <= 16'h0193;    16'd22337: out <= 16'h0409;    16'd22338: out <= 16'hFEE5;    16'd22339: out <= 16'hFFB5;
    16'd22340: out <= 16'h04E4;    16'd22341: out <= 16'h02E2;    16'd22342: out <= 16'h04B3;    16'd22343: out <= 16'h09ED;
    16'd22344: out <= 16'h0345;    16'd22345: out <= 16'h0320;    16'd22346: out <= 16'h0CAA;    16'd22347: out <= 16'h02AF;
    16'd22348: out <= 16'h0132;    16'd22349: out <= 16'h0106;    16'd22350: out <= 16'hFAF1;    16'd22351: out <= 16'h008D;
    16'd22352: out <= 16'hFF23;    16'd22353: out <= 16'h00F2;    16'd22354: out <= 16'h0122;    16'd22355: out <= 16'hFDA0;
    16'd22356: out <= 16'h0803;    16'd22357: out <= 16'h0082;    16'd22358: out <= 16'h0212;    16'd22359: out <= 16'h04DC;
    16'd22360: out <= 16'h084F;    16'd22361: out <= 16'h03AC;    16'd22362: out <= 16'h0442;    16'd22363: out <= 16'h06ED;
    16'd22364: out <= 16'h0657;    16'd22365: out <= 16'h05B8;    16'd22366: out <= 16'h046F;    16'd22367: out <= 16'h0482;
    16'd22368: out <= 16'h040D;    16'd22369: out <= 16'h0413;    16'd22370: out <= 16'h074E;    16'd22371: out <= 16'h02EA;
    16'd22372: out <= 16'h0212;    16'd22373: out <= 16'h05C5;    16'd22374: out <= 16'h01ED;    16'd22375: out <= 16'h0B23;
    16'd22376: out <= 16'h0256;    16'd22377: out <= 16'h0180;    16'd22378: out <= 16'h0376;    16'd22379: out <= 16'h0B40;
    16'd22380: out <= 16'h0972;    16'd22381: out <= 16'h096C;    16'd22382: out <= 16'hFF8B;    16'd22383: out <= 16'h087E;
    16'd22384: out <= 16'h0888;    16'd22385: out <= 16'h05CE;    16'd22386: out <= 16'h02D6;    16'd22387: out <= 16'h04F8;
    16'd22388: out <= 16'h0087;    16'd22389: out <= 16'hFCFA;    16'd22390: out <= 16'hFE6E;    16'd22391: out <= 16'h0C08;
    16'd22392: out <= 16'hFBAF;    16'd22393: out <= 16'h0610;    16'd22394: out <= 16'h046C;    16'd22395: out <= 16'h0C25;
    16'd22396: out <= 16'h0511;    16'd22397: out <= 16'h06DF;    16'd22398: out <= 16'h02D6;    16'd22399: out <= 16'hFE72;
    16'd22400: out <= 16'h090F;    16'd22401: out <= 16'hFF2D;    16'd22402: out <= 16'h02B9;    16'd22403: out <= 16'hFD85;
    16'd22404: out <= 16'h00E9;    16'd22405: out <= 16'h05F6;    16'd22406: out <= 16'h01EC;    16'd22407: out <= 16'h0B84;
    16'd22408: out <= 16'hFF61;    16'd22409: out <= 16'hFD7A;    16'd22410: out <= 16'h05C8;    16'd22411: out <= 16'h0C7F;
    16'd22412: out <= 16'h06A5;    16'd22413: out <= 16'h04AE;    16'd22414: out <= 16'h08B4;    16'd22415: out <= 16'h0565;
    16'd22416: out <= 16'h0A7F;    16'd22417: out <= 16'h0D81;    16'd22418: out <= 16'h0393;    16'd22419: out <= 16'h052F;
    16'd22420: out <= 16'hFAC8;    16'd22421: out <= 16'hFCEA;    16'd22422: out <= 16'h0165;    16'd22423: out <= 16'h030B;
    16'd22424: out <= 16'hFC40;    16'd22425: out <= 16'hF79E;    16'd22426: out <= 16'hFBD5;    16'd22427: out <= 16'h074D;
    16'd22428: out <= 16'h03CE;    16'd22429: out <= 16'h013F;    16'd22430: out <= 16'h02AA;    16'd22431: out <= 16'h012D;
    16'd22432: out <= 16'hFD07;    16'd22433: out <= 16'hFC8D;    16'd22434: out <= 16'h05C0;    16'd22435: out <= 16'h052C;
    16'd22436: out <= 16'hFECB;    16'd22437: out <= 16'h06E7;    16'd22438: out <= 16'h00DF;    16'd22439: out <= 16'h046C;
    16'd22440: out <= 16'hFF26;    16'd22441: out <= 16'h0798;    16'd22442: out <= 16'h00C2;    16'd22443: out <= 16'h0520;
    16'd22444: out <= 16'h03DE;    16'd22445: out <= 16'h08B4;    16'd22446: out <= 16'h0432;    16'd22447: out <= 16'hFF89;
    16'd22448: out <= 16'h064E;    16'd22449: out <= 16'h0443;    16'd22450: out <= 16'h0B53;    16'd22451: out <= 16'h0528;
    16'd22452: out <= 16'h0527;    16'd22453: out <= 16'h0081;    16'd22454: out <= 16'h0401;    16'd22455: out <= 16'h099C;
    16'd22456: out <= 16'h0343;    16'd22457: out <= 16'h07AF;    16'd22458: out <= 16'h0408;    16'd22459: out <= 16'h06B6;
    16'd22460: out <= 16'hFDDA;    16'd22461: out <= 16'h069B;    16'd22462: out <= 16'h07F4;    16'd22463: out <= 16'h028A;
    16'd22464: out <= 16'h06D9;    16'd22465: out <= 16'h0161;    16'd22466: out <= 16'h0520;    16'd22467: out <= 16'h03E9;
    16'd22468: out <= 16'h0619;    16'd22469: out <= 16'hFF9D;    16'd22470: out <= 16'h0353;    16'd22471: out <= 16'h0306;
    16'd22472: out <= 16'h01BE;    16'd22473: out <= 16'h0540;    16'd22474: out <= 16'h018C;    16'd22475: out <= 16'h00E4;
    16'd22476: out <= 16'h0580;    16'd22477: out <= 16'h05A9;    16'd22478: out <= 16'h054C;    16'd22479: out <= 16'h03F9;
    16'd22480: out <= 16'hF9EA;    16'd22481: out <= 16'h0768;    16'd22482: out <= 16'h030B;    16'd22483: out <= 16'h0460;
    16'd22484: out <= 16'h0169;    16'd22485: out <= 16'h05CF;    16'd22486: out <= 16'h0430;    16'd22487: out <= 16'h059D;
    16'd22488: out <= 16'hFB83;    16'd22489: out <= 16'hFDBD;    16'd22490: out <= 16'hFFAE;    16'd22491: out <= 16'hF7B6;
    16'd22492: out <= 16'hFC12;    16'd22493: out <= 16'hF7E8;    16'd22494: out <= 16'hFCAB;    16'd22495: out <= 16'h042D;
    16'd22496: out <= 16'hFF11;    16'd22497: out <= 16'h0463;    16'd22498: out <= 16'h01C6;    16'd22499: out <= 16'h00F1;
    16'd22500: out <= 16'hFF24;    16'd22501: out <= 16'hFCD1;    16'd22502: out <= 16'h0041;    16'd22503: out <= 16'h0064;
    16'd22504: out <= 16'h04E1;    16'd22505: out <= 16'h03BA;    16'd22506: out <= 16'h006B;    16'd22507: out <= 16'hFD24;
    16'd22508: out <= 16'h01ED;    16'd22509: out <= 16'hFC3F;    16'd22510: out <= 16'h0364;    16'd22511: out <= 16'h0533;
    16'd22512: out <= 16'h02AF;    16'd22513: out <= 16'hFBC3;    16'd22514: out <= 16'h00D9;    16'd22515: out <= 16'h079F;
    16'd22516: out <= 16'hF934;    16'd22517: out <= 16'hFB90;    16'd22518: out <= 16'h042A;    16'd22519: out <= 16'h0329;
    16'd22520: out <= 16'h023D;    16'd22521: out <= 16'hFD67;    16'd22522: out <= 16'hFE70;    16'd22523: out <= 16'hFFDC;
    16'd22524: out <= 16'hFD21;    16'd22525: out <= 16'h05A7;    16'd22526: out <= 16'h02DF;    16'd22527: out <= 16'h049B;
    16'd22528: out <= 16'h00F8;    16'd22529: out <= 16'h0892;    16'd22530: out <= 16'hF75F;    16'd22531: out <= 16'h018F;
    16'd22532: out <= 16'hF4CA;    16'd22533: out <= 16'h0011;    16'd22534: out <= 16'hFB9D;    16'd22535: out <= 16'hFFB0;
    16'd22536: out <= 16'hFDC0;    16'd22537: out <= 16'hFC37;    16'd22538: out <= 16'hFE5E;    16'd22539: out <= 16'h023F;
    16'd22540: out <= 16'hFBEA;    16'd22541: out <= 16'h080F;    16'd22542: out <= 16'h018E;    16'd22543: out <= 16'h00ED;
    16'd22544: out <= 16'h01C3;    16'd22545: out <= 16'h0119;    16'd22546: out <= 16'hF8AF;    16'd22547: out <= 16'h00F7;
    16'd22548: out <= 16'h04A4;    16'd22549: out <= 16'h039B;    16'd22550: out <= 16'hFDA9;    16'd22551: out <= 16'hFDA4;
    16'd22552: out <= 16'h026D;    16'd22553: out <= 16'h0292;    16'd22554: out <= 16'h02AC;    16'd22555: out <= 16'hFDBC;
    16'd22556: out <= 16'hFD88;    16'd22557: out <= 16'h0146;    16'd22558: out <= 16'h0394;    16'd22559: out <= 16'h0328;
    16'd22560: out <= 16'h01D3;    16'd22561: out <= 16'h069B;    16'd22562: out <= 16'h02EC;    16'd22563: out <= 16'h06F8;
    16'd22564: out <= 16'h08AD;    16'd22565: out <= 16'h03E1;    16'd22566: out <= 16'h0197;    16'd22567: out <= 16'h05E1;
    16'd22568: out <= 16'hFD42;    16'd22569: out <= 16'h0CFF;    16'd22570: out <= 16'h02E5;    16'd22571: out <= 16'h0900;
    16'd22572: out <= 16'h090C;    16'd22573: out <= 16'h0317;    16'd22574: out <= 16'h0994;    16'd22575: out <= 16'h040A;
    16'd22576: out <= 16'h07D8;    16'd22577: out <= 16'h0742;    16'd22578: out <= 16'h027B;    16'd22579: out <= 16'hFFDF;
    16'd22580: out <= 16'h0645;    16'd22581: out <= 16'h0322;    16'd22582: out <= 16'h010E;    16'd22583: out <= 16'hFFB4;
    16'd22584: out <= 16'h0634;    16'd22585: out <= 16'h06CC;    16'd22586: out <= 16'h010F;    16'd22587: out <= 16'hFF37;
    16'd22588: out <= 16'h067D;    16'd22589: out <= 16'h0005;    16'd22590: out <= 16'h05F9;    16'd22591: out <= 16'h0509;
    16'd22592: out <= 16'h0411;    16'd22593: out <= 16'h0738;    16'd22594: out <= 16'h025E;    16'd22595: out <= 16'h062C;
    16'd22596: out <= 16'h0901;    16'd22597: out <= 16'h0420;    16'd22598: out <= 16'hFCB3;    16'd22599: out <= 16'h02E1;
    16'd22600: out <= 16'h0315;    16'd22601: out <= 16'hFD9F;    16'd22602: out <= 16'h036A;    16'd22603: out <= 16'h08AC;
    16'd22604: out <= 16'h0397;    16'd22605: out <= 16'h0539;    16'd22606: out <= 16'h02FB;    16'd22607: out <= 16'hF994;
    16'd22608: out <= 16'h0012;    16'd22609: out <= 16'h034E;    16'd22610: out <= 16'h0691;    16'd22611: out <= 16'hFFA1;
    16'd22612: out <= 16'h0391;    16'd22613: out <= 16'h06E7;    16'd22614: out <= 16'h05FD;    16'd22615: out <= 16'h02C3;
    16'd22616: out <= 16'h06DD;    16'd22617: out <= 16'h075D;    16'd22618: out <= 16'h01C8;    16'd22619: out <= 16'h0939;
    16'd22620: out <= 16'hFF05;    16'd22621: out <= 16'hFDBF;    16'd22622: out <= 16'h056B;    16'd22623: out <= 16'h0851;
    16'd22624: out <= 16'h02D7;    16'd22625: out <= 16'h0025;    16'd22626: out <= 16'h031B;    16'd22627: out <= 16'hFFA1;
    16'd22628: out <= 16'h01E6;    16'd22629: out <= 16'hFBAF;    16'd22630: out <= 16'hFB92;    16'd22631: out <= 16'h002B;
    16'd22632: out <= 16'h02B3;    16'd22633: out <= 16'h03E6;    16'd22634: out <= 16'hFED0;    16'd22635: out <= 16'h0392;
    16'd22636: out <= 16'h0385;    16'd22637: out <= 16'h0295;    16'd22638: out <= 16'h1159;    16'd22639: out <= 16'h03ED;
    16'd22640: out <= 16'h023B;    16'd22641: out <= 16'h0A42;    16'd22642: out <= 16'h0712;    16'd22643: out <= 16'h06CA;
    16'd22644: out <= 16'hFB3E;    16'd22645: out <= 16'h070A;    16'd22646: out <= 16'h05C5;    16'd22647: out <= 16'h050A;
    16'd22648: out <= 16'h0740;    16'd22649: out <= 16'hFC8B;    16'd22650: out <= 16'h0324;    16'd22651: out <= 16'h0138;
    16'd22652: out <= 16'h038E;    16'd22653: out <= 16'h05CE;    16'd22654: out <= 16'h0135;    16'd22655: out <= 16'h0153;
    16'd22656: out <= 16'h0350;    16'd22657: out <= 16'h0503;    16'd22658: out <= 16'h0261;    16'd22659: out <= 16'h0354;
    16'd22660: out <= 16'h061D;    16'd22661: out <= 16'h00FD;    16'd22662: out <= 16'h0532;    16'd22663: out <= 16'h0080;
    16'd22664: out <= 16'hFDA0;    16'd22665: out <= 16'hFFCD;    16'd22666: out <= 16'hFFB7;    16'd22667: out <= 16'h044D;
    16'd22668: out <= 16'h069E;    16'd22669: out <= 16'h082B;    16'd22670: out <= 16'h0798;    16'd22671: out <= 16'h082D;
    16'd22672: out <= 16'h006B;    16'd22673: out <= 16'hFFF5;    16'd22674: out <= 16'hFAAD;    16'd22675: out <= 16'h056F;
    16'd22676: out <= 16'hFCD1;    16'd22677: out <= 16'h03F8;    16'd22678: out <= 16'hFE47;    16'd22679: out <= 16'hFE6C;
    16'd22680: out <= 16'hFDCA;    16'd22681: out <= 16'h00D4;    16'd22682: out <= 16'hFF5F;    16'd22683: out <= 16'h0108;
    16'd22684: out <= 16'h0060;    16'd22685: out <= 16'h049D;    16'd22686: out <= 16'hFCC9;    16'd22687: out <= 16'hFF70;
    16'd22688: out <= 16'h026A;    16'd22689: out <= 16'h01A2;    16'd22690: out <= 16'h0367;    16'd22691: out <= 16'hFEF3;
    16'd22692: out <= 16'hFD31;    16'd22693: out <= 16'h0289;    16'd22694: out <= 16'hFA24;    16'd22695: out <= 16'hFB8C;
    16'd22696: out <= 16'hFC68;    16'd22697: out <= 16'h00C0;    16'd22698: out <= 16'h039C;    16'd22699: out <= 16'h02FD;
    16'd22700: out <= 16'hFD9A;    16'd22701: out <= 16'h000B;    16'd22702: out <= 16'hFDE3;    16'd22703: out <= 16'h0280;
    16'd22704: out <= 16'h07DB;    16'd22705: out <= 16'h0012;    16'd22706: out <= 16'h00B8;    16'd22707: out <= 16'h075E;
    16'd22708: out <= 16'h02BA;    16'd22709: out <= 16'h0411;    16'd22710: out <= 16'h05ED;    16'd22711: out <= 16'h0353;
    16'd22712: out <= 16'h0475;    16'd22713: out <= 16'h05EA;    16'd22714: out <= 16'h04A1;    16'd22715: out <= 16'h0315;
    16'd22716: out <= 16'h0765;    16'd22717: out <= 16'h046A;    16'd22718: out <= 16'h01B4;    16'd22719: out <= 16'hFFAC;
    16'd22720: out <= 16'h0E72;    16'd22721: out <= 16'h014C;    16'd22722: out <= 16'h0B60;    16'd22723: out <= 16'h01D2;
    16'd22724: out <= 16'h024D;    16'd22725: out <= 16'h039F;    16'd22726: out <= 16'h0155;    16'd22727: out <= 16'h0B5F;
    16'd22728: out <= 16'h0669;    16'd22729: out <= 16'h06A4;    16'd22730: out <= 16'h0288;    16'd22731: out <= 16'h04EA;
    16'd22732: out <= 16'h047B;    16'd22733: out <= 16'hF9E9;    16'd22734: out <= 16'h030F;    16'd22735: out <= 16'h0918;
    16'd22736: out <= 16'h097F;    16'd22737: out <= 16'h05DC;    16'd22738: out <= 16'hFCF1;    16'd22739: out <= 16'h0345;
    16'd22740: out <= 16'hFF3A;    16'd22741: out <= 16'h07C4;    16'd22742: out <= 16'h08DC;    16'd22743: out <= 16'h0274;
    16'd22744: out <= 16'h060B;    16'd22745: out <= 16'h0454;    16'd22746: out <= 16'hFE14;    16'd22747: out <= 16'hFB42;
    16'd22748: out <= 16'hFE53;    16'd22749: out <= 16'h02C6;    16'd22750: out <= 16'h02C0;    16'd22751: out <= 16'hFCBF;
    16'd22752: out <= 16'hFE05;    16'd22753: out <= 16'h027B;    16'd22754: out <= 16'h0465;    16'd22755: out <= 16'h0011;
    16'd22756: out <= 16'h0438;    16'd22757: out <= 16'h00FB;    16'd22758: out <= 16'hFD5C;    16'd22759: out <= 16'h04C5;
    16'd22760: out <= 16'h0107;    16'd22761: out <= 16'h02C1;    16'd22762: out <= 16'hFF58;    16'd22763: out <= 16'h02C0;
    16'd22764: out <= 16'hFAAB;    16'd22765: out <= 16'hF91F;    16'd22766: out <= 16'hFBC6;    16'd22767: out <= 16'h0088;
    16'd22768: out <= 16'h00C4;    16'd22769: out <= 16'h0222;    16'd22770: out <= 16'hFCE3;    16'd22771: out <= 16'hFC7E;
    16'd22772: out <= 16'h05DC;    16'd22773: out <= 16'hF964;    16'd22774: out <= 16'hFE4B;    16'd22775: out <= 16'h01D3;
    16'd22776: out <= 16'h02B2;    16'd22777: out <= 16'h0568;    16'd22778: out <= 16'hFE8D;    16'd22779: out <= 16'h0646;
    16'd22780: out <= 16'h00AE;    16'd22781: out <= 16'hFAB6;    16'd22782: out <= 16'hFF06;    16'd22783: out <= 16'hFE77;
    16'd22784: out <= 16'h0455;    16'd22785: out <= 16'h0217;    16'd22786: out <= 16'h06B1;    16'd22787: out <= 16'hFD33;
    16'd22788: out <= 16'hFC7C;    16'd22789: out <= 16'h0414;    16'd22790: out <= 16'hFF57;    16'd22791: out <= 16'h0170;
    16'd22792: out <= 16'h02AD;    16'd22793: out <= 16'hFF75;    16'd22794: out <= 16'hF7C5;    16'd22795: out <= 16'h0326;
    16'd22796: out <= 16'h06F2;    16'd22797: out <= 16'h073A;    16'd22798: out <= 16'hF9E0;    16'd22799: out <= 16'h0214;
    16'd22800: out <= 16'h01E3;    16'd22801: out <= 16'h03D7;    16'd22802: out <= 16'h04F4;    16'd22803: out <= 16'h029F;
    16'd22804: out <= 16'hFDC4;    16'd22805: out <= 16'hFA66;    16'd22806: out <= 16'h02F4;    16'd22807: out <= 16'hFF77;
    16'd22808: out <= 16'hFFBF;    16'd22809: out <= 16'h008F;    16'd22810: out <= 16'hFA3B;    16'd22811: out <= 16'h001A;
    16'd22812: out <= 16'h0B45;    16'd22813: out <= 16'h10D2;    16'd22814: out <= 16'h0B95;    16'd22815: out <= 16'h0827;
    16'd22816: out <= 16'h0685;    16'd22817: out <= 16'h0C73;    16'd22818: out <= 16'h09F9;    16'd22819: out <= 16'h0D50;
    16'd22820: out <= 16'h05C1;    16'd22821: out <= 16'h055D;    16'd22822: out <= 16'h04C9;    16'd22823: out <= 16'h032A;
    16'd22824: out <= 16'hFFA6;    16'd22825: out <= 16'h03F9;    16'd22826: out <= 16'h00BF;    16'd22827: out <= 16'h0714;
    16'd22828: out <= 16'h085E;    16'd22829: out <= 16'h047A;    16'd22830: out <= 16'h072C;    16'd22831: out <= 16'h0277;
    16'd22832: out <= 16'h0657;    16'd22833: out <= 16'h0A7E;    16'd22834: out <= 16'h051C;    16'd22835: out <= 16'h0468;
    16'd22836: out <= 16'h046D;    16'd22837: out <= 16'h0332;    16'd22838: out <= 16'h06C0;    16'd22839: out <= 16'h020F;
    16'd22840: out <= 16'hFBCF;    16'd22841: out <= 16'h0460;    16'd22842: out <= 16'h0834;    16'd22843: out <= 16'h03DE;
    16'd22844: out <= 16'hFFA1;    16'd22845: out <= 16'h0244;    16'd22846: out <= 16'h0623;    16'd22847: out <= 16'h0D6A;
    16'd22848: out <= 16'h067D;    16'd22849: out <= 16'h04C2;    16'd22850: out <= 16'h0A28;    16'd22851: out <= 16'h0291;
    16'd22852: out <= 16'hFEE2;    16'd22853: out <= 16'h06FB;    16'd22854: out <= 16'h021C;    16'd22855: out <= 16'h09B1;
    16'd22856: out <= 16'h0397;    16'd22857: out <= 16'h0569;    16'd22858: out <= 16'hFE1B;    16'd22859: out <= 16'h0278;
    16'd22860: out <= 16'h014F;    16'd22861: out <= 16'h03F4;    16'd22862: out <= 16'hFEA4;    16'd22863: out <= 16'h09BA;
    16'd22864: out <= 16'hFFC1;    16'd22865: out <= 16'h0BCE;    16'd22866: out <= 16'h083C;    16'd22867: out <= 16'h0279;
    16'd22868: out <= 16'hFCB7;    16'd22869: out <= 16'h08C5;    16'd22870: out <= 16'h0C83;    16'd22871: out <= 16'h041A;
    16'd22872: out <= 16'h0308;    16'd22873: out <= 16'h0719;    16'd22874: out <= 16'h05AA;    16'd22875: out <= 16'hFD9A;
    16'd22876: out <= 16'hFE99;    16'd22877: out <= 16'hFE98;    16'd22878: out <= 16'h0B9A;    16'd22879: out <= 16'hFFBB;
    16'd22880: out <= 16'h0355;    16'd22881: out <= 16'h046E;    16'd22882: out <= 16'h0812;    16'd22883: out <= 16'hFFA1;
    16'd22884: out <= 16'h00F1;    16'd22885: out <= 16'h0795;    16'd22886: out <= 16'h004D;    16'd22887: out <= 16'h009A;
    16'd22888: out <= 16'hFE4F;    16'd22889: out <= 16'h05E3;    16'd22890: out <= 16'h0715;    16'd22891: out <= 16'h0A7C;
    16'd22892: out <= 16'h0541;    16'd22893: out <= 16'h061A;    16'd22894: out <= 16'hFACF;    16'd22895: out <= 16'h0259;
    16'd22896: out <= 16'h0965;    16'd22897: out <= 16'h0552;    16'd22898: out <= 16'hFDB3;    16'd22899: out <= 16'h04FC;
    16'd22900: out <= 16'h0019;    16'd22901: out <= 16'h018C;    16'd22902: out <= 16'hFFB6;    16'd22903: out <= 16'hFF79;
    16'd22904: out <= 16'h04A6;    16'd22905: out <= 16'hFD73;    16'd22906: out <= 16'h06BA;    16'd22907: out <= 16'h03D5;
    16'd22908: out <= 16'h0385;    16'd22909: out <= 16'h040E;    16'd22910: out <= 16'h0127;    16'd22911: out <= 16'h014A;
    16'd22912: out <= 16'h02DE;    16'd22913: out <= 16'h0270;    16'd22914: out <= 16'h0232;    16'd22915: out <= 16'h0678;
    16'd22916: out <= 16'h0600;    16'd22917: out <= 16'h042C;    16'd22918: out <= 16'h00B2;    16'd22919: out <= 16'hFAC8;
    16'd22920: out <= 16'h0B64;    16'd22921: out <= 16'h089F;    16'd22922: out <= 16'h0229;    16'd22923: out <= 16'h0165;
    16'd22924: out <= 16'h02D9;    16'd22925: out <= 16'h027D;    16'd22926: out <= 16'hFD84;    16'd22927: out <= 16'h00D7;
    16'd22928: out <= 16'h06F2;    16'd22929: out <= 16'h037A;    16'd22930: out <= 16'h0066;    16'd22931: out <= 16'hFF94;
    16'd22932: out <= 16'h027E;    16'd22933: out <= 16'hF95D;    16'd22934: out <= 16'h006A;    16'd22935: out <= 16'hFF77;
    16'd22936: out <= 16'h014E;    16'd22937: out <= 16'hF6C9;    16'd22938: out <= 16'h0040;    16'd22939: out <= 16'h021D;
    16'd22940: out <= 16'h0879;    16'd22941: out <= 16'h069E;    16'd22942: out <= 16'hFD36;    16'd22943: out <= 16'hFD16;
    16'd22944: out <= 16'hFD24;    16'd22945: out <= 16'h00AE;    16'd22946: out <= 16'h028C;    16'd22947: out <= 16'h05FE;
    16'd22948: out <= 16'h0213;    16'd22949: out <= 16'hFF2B;    16'd22950: out <= 16'h044D;    16'd22951: out <= 16'h0C1B;
    16'd22952: out <= 16'h0A43;    16'd22953: out <= 16'h0858;    16'd22954: out <= 16'h07F8;    16'd22955: out <= 16'h0056;
    16'd22956: out <= 16'h00C7;    16'd22957: out <= 16'h007B;    16'd22958: out <= 16'h062A;    16'd22959: out <= 16'h06C0;
    16'd22960: out <= 16'h0260;    16'd22961: out <= 16'h0095;    16'd22962: out <= 16'h0B4D;    16'd22963: out <= 16'h01CC;
    16'd22964: out <= 16'hFC22;    16'd22965: out <= 16'h09F5;    16'd22966: out <= 16'h032A;    16'd22967: out <= 16'h0704;
    16'd22968: out <= 16'h088C;    16'd22969: out <= 16'h0239;    16'd22970: out <= 16'h0863;    16'd22971: out <= 16'h0734;
    16'd22972: out <= 16'h0B22;    16'd22973: out <= 16'h00F1;    16'd22974: out <= 16'h0B2C;    16'd22975: out <= 16'h029F;
    16'd22976: out <= 16'hFFB2;    16'd22977: out <= 16'h07C1;    16'd22978: out <= 16'h0291;    16'd22979: out <= 16'h0A57;
    16'd22980: out <= 16'h07F5;    16'd22981: out <= 16'h0AF1;    16'd22982: out <= 16'h0088;    16'd22983: out <= 16'h046B;
    16'd22984: out <= 16'h03F4;    16'd22985: out <= 16'h0615;    16'd22986: out <= 16'h0476;    16'd22987: out <= 16'h0690;
    16'd22988: out <= 16'h00FC;    16'd22989: out <= 16'h0976;    16'd22990: out <= 16'h05D3;    16'd22991: out <= 16'h07DB;
    16'd22992: out <= 16'h079A;    16'd22993: out <= 16'h0283;    16'd22994: out <= 16'hFFE8;    16'd22995: out <= 16'h0613;
    16'd22996: out <= 16'h0897;    16'd22997: out <= 16'hFDD2;    16'd22998: out <= 16'h0454;    16'd22999: out <= 16'h03B5;
    16'd23000: out <= 16'h09B8;    16'd23001: out <= 16'h0111;    16'd23002: out <= 16'h0720;    16'd23003: out <= 16'h01AE;
    16'd23004: out <= 16'hFE9A;    16'd23005: out <= 16'hFF0E;    16'd23006: out <= 16'h0415;    16'd23007: out <= 16'hFD0A;
    16'd23008: out <= 16'hFC5A;    16'd23009: out <= 16'hFD8B;    16'd23010: out <= 16'h0088;    16'd23011: out <= 16'hFA1A;
    16'd23012: out <= 16'h0370;    16'd23013: out <= 16'hFD8A;    16'd23014: out <= 16'h03CB;    16'd23015: out <= 16'hFCE0;
    16'd23016: out <= 16'h012F;    16'd23017: out <= 16'hFF0D;    16'd23018: out <= 16'h0080;    16'd23019: out <= 16'hFF20;
    16'd23020: out <= 16'h01F2;    16'd23021: out <= 16'h040A;    16'd23022: out <= 16'hFFB8;    16'd23023: out <= 16'hFD62;
    16'd23024: out <= 16'hFD8B;    16'd23025: out <= 16'hFE93;    16'd23026: out <= 16'h01E1;    16'd23027: out <= 16'hFCDE;
    16'd23028: out <= 16'hFDDB;    16'd23029: out <= 16'h0296;    16'd23030: out <= 16'hFCB9;    16'd23031: out <= 16'h0318;
    16'd23032: out <= 16'h01ED;    16'd23033: out <= 16'hFE05;    16'd23034: out <= 16'h01FD;    16'd23035: out <= 16'hF92A;
    16'd23036: out <= 16'h0366;    16'd23037: out <= 16'h007E;    16'd23038: out <= 16'hFF24;    16'd23039: out <= 16'h024E;
    16'd23040: out <= 16'h07DD;    16'd23041: out <= 16'h0672;    16'd23042: out <= 16'hFBC9;    16'd23043: out <= 16'hFF14;
    16'd23044: out <= 16'h0818;    16'd23045: out <= 16'h0211;    16'd23046: out <= 16'h0058;    16'd23047: out <= 16'hFCBD;
    16'd23048: out <= 16'hFFFA;    16'd23049: out <= 16'hFE18;    16'd23050: out <= 16'h03CF;    16'd23051: out <= 16'hFB4A;
    16'd23052: out <= 16'hFF5B;    16'd23053: out <= 16'h0217;    16'd23054: out <= 16'h0412;    16'd23055: out <= 16'h01AC;
    16'd23056: out <= 16'hFE5E;    16'd23057: out <= 16'hFC2E;    16'd23058: out <= 16'h051D;    16'd23059: out <= 16'h020F;
    16'd23060: out <= 16'h07D2;    16'd23061: out <= 16'h01E8;    16'd23062: out <= 16'hF8D0;    16'd23063: out <= 16'hF9D6;
    16'd23064: out <= 16'h010A;    16'd23065: out <= 16'h00EC;    16'd23066: out <= 16'h0069;    16'd23067: out <= 16'h0764;
    16'd23068: out <= 16'h021A;    16'd23069: out <= 16'h08CF;    16'd23070: out <= 16'h05B6;    16'd23071: out <= 16'h0CEA;
    16'd23072: out <= 16'h02F2;    16'd23073: out <= 16'h0167;    16'd23074: out <= 16'h04E8;    16'd23075: out <= 16'h02F7;
    16'd23076: out <= 16'h0237;    16'd23077: out <= 16'h001F;    16'd23078: out <= 16'h09ED;    16'd23079: out <= 16'h03EB;
    16'd23080: out <= 16'h0498;    16'd23081: out <= 16'h0353;    16'd23082: out <= 16'h06E3;    16'd23083: out <= 16'h08B8;
    16'd23084: out <= 16'h08B8;    16'd23085: out <= 16'h02B1;    16'd23086: out <= 16'h0156;    16'd23087: out <= 16'h0498;
    16'd23088: out <= 16'h06F4;    16'd23089: out <= 16'h0586;    16'd23090: out <= 16'h0355;    16'd23091: out <= 16'h0472;
    16'd23092: out <= 16'h07E6;    16'd23093: out <= 16'h06FE;    16'd23094: out <= 16'h0638;    16'd23095: out <= 16'hFF1B;
    16'd23096: out <= 16'hFE98;    16'd23097: out <= 16'h07DB;    16'd23098: out <= 16'hFB6C;    16'd23099: out <= 16'h02D1;
    16'd23100: out <= 16'h06AF;    16'd23101: out <= 16'h07D5;    16'd23102: out <= 16'h0291;    16'd23103: out <= 16'h067B;
    16'd23104: out <= 16'h0511;    16'd23105: out <= 16'h0988;    16'd23106: out <= 16'h0519;    16'd23107: out <= 16'h049D;
    16'd23108: out <= 16'h06CE;    16'd23109: out <= 16'h0393;    16'd23110: out <= 16'h0AED;    16'd23111: out <= 16'h0463;
    16'd23112: out <= 16'hFFAA;    16'd23113: out <= 16'h05DD;    16'd23114: out <= 16'h01D4;    16'd23115: out <= 16'h02E8;
    16'd23116: out <= 16'h048A;    16'd23117: out <= 16'h0575;    16'd23118: out <= 16'h058E;    16'd23119: out <= 16'h008B;
    16'd23120: out <= 16'h005D;    16'd23121: out <= 16'h0356;    16'd23122: out <= 16'h07CB;    16'd23123: out <= 16'h074D;
    16'd23124: out <= 16'h0916;    16'd23125: out <= 16'h023D;    16'd23126: out <= 16'h027B;    16'd23127: out <= 16'h01C7;
    16'd23128: out <= 16'h0A5C;    16'd23129: out <= 16'h0414;    16'd23130: out <= 16'hFEA6;    16'd23131: out <= 16'h0477;
    16'd23132: out <= 16'h08C4;    16'd23133: out <= 16'hFFB9;    16'd23134: out <= 16'h07F1;    16'd23135: out <= 16'h0010;
    16'd23136: out <= 16'h0705;    16'd23137: out <= 16'h001F;    16'd23138: out <= 16'h0993;    16'd23139: out <= 16'hFF14;
    16'd23140: out <= 16'h0715;    16'd23141: out <= 16'h0A59;    16'd23142: out <= 16'h0478;    16'd23143: out <= 16'h000D;
    16'd23144: out <= 16'h01DF;    16'd23145: out <= 16'h064D;    16'd23146: out <= 16'h06A0;    16'd23147: out <= 16'hFE9B;
    16'd23148: out <= 16'h05FD;    16'd23149: out <= 16'hFED1;    16'd23150: out <= 16'h0650;    16'd23151: out <= 16'h0045;
    16'd23152: out <= 16'h0434;    16'd23153: out <= 16'hFCEE;    16'd23154: out <= 16'h0426;    16'd23155: out <= 16'hFDE1;
    16'd23156: out <= 16'h016E;    16'd23157: out <= 16'h0234;    16'd23158: out <= 16'h023B;    16'd23159: out <= 16'h054F;
    16'd23160: out <= 16'h00AF;    16'd23161: out <= 16'h0778;    16'd23162: out <= 16'h043F;    16'd23163: out <= 16'h0761;
    16'd23164: out <= 16'h05B8;    16'd23165: out <= 16'h027A;    16'd23166: out <= 16'h0170;    16'd23167: out <= 16'h07DF;
    16'd23168: out <= 16'h0670;    16'd23169: out <= 16'h00F4;    16'd23170: out <= 16'h030D;    16'd23171: out <= 16'h01EE;
    16'd23172: out <= 16'h0271;    16'd23173: out <= 16'h0990;    16'd23174: out <= 16'h0443;    16'd23175: out <= 16'h03A6;
    16'd23176: out <= 16'hFB16;    16'd23177: out <= 16'hFFD1;    16'd23178: out <= 16'h03EE;    16'd23179: out <= 16'h000D;
    16'd23180: out <= 16'h04A2;    16'd23181: out <= 16'h0492;    16'd23182: out <= 16'h0B7A;    16'd23183: out <= 16'h0A92;
    16'd23184: out <= 16'h0117;    16'd23185: out <= 16'h0870;    16'd23186: out <= 16'h0115;    16'd23187: out <= 16'h009B;
    16'd23188: out <= 16'hFF6C;    16'd23189: out <= 16'h0067;    16'd23190: out <= 16'h0081;    16'd23191: out <= 16'hFC71;
    16'd23192: out <= 16'hFEF2;    16'd23193: out <= 16'hFF8A;    16'd23194: out <= 16'h0B5C;    16'd23195: out <= 16'hFC3B;
    16'd23196: out <= 16'hF998;    16'd23197: out <= 16'h0445;    16'd23198: out <= 16'h0267;    16'd23199: out <= 16'h0340;
    16'd23200: out <= 16'hFE39;    16'd23201: out <= 16'hFEE7;    16'd23202: out <= 16'h0091;    16'd23203: out <= 16'h03B6;
    16'd23204: out <= 16'h03B7;    16'd23205: out <= 16'h0487;    16'd23206: out <= 16'h0061;    16'd23207: out <= 16'h055C;
    16'd23208: out <= 16'h05ED;    16'd23209: out <= 16'h051F;    16'd23210: out <= 16'h0724;    16'd23211: out <= 16'h06A1;
    16'd23212: out <= 16'h0534;    16'd23213: out <= 16'h01B4;    16'd23214: out <= 16'h01FD;    16'd23215: out <= 16'h03BD;
    16'd23216: out <= 16'h007A;    16'd23217: out <= 16'h048C;    16'd23218: out <= 16'h04FF;    16'd23219: out <= 16'h0669;
    16'd23220: out <= 16'h06E4;    16'd23221: out <= 16'h0A72;    16'd23222: out <= 16'h09C4;    16'd23223: out <= 16'h05BF;
    16'd23224: out <= 16'hFFAA;    16'd23225: out <= 16'h0084;    16'd23226: out <= 16'h0384;    16'd23227: out <= 16'h0595;
    16'd23228: out <= 16'h06F6;    16'd23229: out <= 16'h04E7;    16'd23230: out <= 16'h07F6;    16'd23231: out <= 16'h0325;
    16'd23232: out <= 16'h04E6;    16'd23233: out <= 16'h05C1;    16'd23234: out <= 16'h0517;    16'd23235: out <= 16'h0908;
    16'd23236: out <= 16'h04D9;    16'd23237: out <= 16'h07A9;    16'd23238: out <= 16'hFE0D;    16'd23239: out <= 16'h04D4;
    16'd23240: out <= 16'h052F;    16'd23241: out <= 16'hFE0C;    16'd23242: out <= 16'hFE89;    16'd23243: out <= 16'h05E1;
    16'd23244: out <= 16'h0753;    16'd23245: out <= 16'h050D;    16'd23246: out <= 16'h07ED;    16'd23247: out <= 16'h0666;
    16'd23248: out <= 16'h0736;    16'd23249: out <= 16'h0169;    16'd23250: out <= 16'h033F;    16'd23251: out <= 16'hFDBA;
    16'd23252: out <= 16'h06F4;    16'd23253: out <= 16'hFCDC;    16'd23254: out <= 16'hFA66;    16'd23255: out <= 16'h00F9;
    16'd23256: out <= 16'h03F9;    16'd23257: out <= 16'hFE59;    16'd23258: out <= 16'h0273;    16'd23259: out <= 16'h0093;
    16'd23260: out <= 16'hFFD9;    16'd23261: out <= 16'hFB1F;    16'd23262: out <= 16'hFE01;    16'd23263: out <= 16'h045F;
    16'd23264: out <= 16'hFAA3;    16'd23265: out <= 16'h0271;    16'd23266: out <= 16'h00E9;    16'd23267: out <= 16'h0482;
    16'd23268: out <= 16'h05FB;    16'd23269: out <= 16'hFE36;    16'd23270: out <= 16'h06C8;    16'd23271: out <= 16'h06AC;
    16'd23272: out <= 16'h0595;    16'd23273: out <= 16'h05C3;    16'd23274: out <= 16'hFDE5;    16'd23275: out <= 16'h0766;
    16'd23276: out <= 16'hFE15;    16'd23277: out <= 16'hFB0F;    16'd23278: out <= 16'hFEA4;    16'd23279: out <= 16'hFBD4;
    16'd23280: out <= 16'h0737;    16'd23281: out <= 16'hF704;    16'd23282: out <= 16'hFFF7;    16'd23283: out <= 16'hFB3F;
    16'd23284: out <= 16'hFEFE;    16'd23285: out <= 16'hF82C;    16'd23286: out <= 16'h05B6;    16'd23287: out <= 16'hFBEE;
    16'd23288: out <= 16'hFF49;    16'd23289: out <= 16'hFB47;    16'd23290: out <= 16'hFF80;    16'd23291: out <= 16'hFFFB;
    16'd23292: out <= 16'h0151;    16'd23293: out <= 16'h0028;    16'd23294: out <= 16'hFBCD;    16'd23295: out <= 16'h0015;
    16'd23296: out <= 16'h00A5;    16'd23297: out <= 16'h023C;    16'd23298: out <= 16'h0246;    16'd23299: out <= 16'h032A;
    16'd23300: out <= 16'hFE71;    16'd23301: out <= 16'hFCCE;    16'd23302: out <= 16'hFD42;    16'd23303: out <= 16'hF937;
    16'd23304: out <= 16'h00E9;    16'd23305: out <= 16'h04BA;    16'd23306: out <= 16'hFD11;    16'd23307: out <= 16'hFDA7;
    16'd23308: out <= 16'h0569;    16'd23309: out <= 16'h0297;    16'd23310: out <= 16'h070D;    16'd23311: out <= 16'h028B;
    16'd23312: out <= 16'hFBC4;    16'd23313: out <= 16'hFA8C;    16'd23314: out <= 16'hFED4;    16'd23315: out <= 16'h021E;
    16'd23316: out <= 16'hFF8E;    16'd23317: out <= 16'hF770;    16'd23318: out <= 16'h03D7;    16'd23319: out <= 16'h0645;
    16'd23320: out <= 16'h01A0;    16'd23321: out <= 16'h032C;    16'd23322: out <= 16'h0542;    16'd23323: out <= 16'h0244;
    16'd23324: out <= 16'h00C8;    16'd23325: out <= 16'hFD9E;    16'd23326: out <= 16'h0711;    16'd23327: out <= 16'hFDC2;
    16'd23328: out <= 16'h05FE;    16'd23329: out <= 16'h0605;    16'd23330: out <= 16'hFEF4;    16'd23331: out <= 16'hFCC1;
    16'd23332: out <= 16'h0773;    16'd23333: out <= 16'h042B;    16'd23334: out <= 16'h013D;    16'd23335: out <= 16'h09E5;
    16'd23336: out <= 16'h03F4;    16'd23337: out <= 16'h012F;    16'd23338: out <= 16'h0471;    16'd23339: out <= 16'h02B9;
    16'd23340: out <= 16'h04C1;    16'd23341: out <= 16'h00E9;    16'd23342: out <= 16'h056B;    16'd23343: out <= 16'h05C7;
    16'd23344: out <= 16'h09CF;    16'd23345: out <= 16'h09DE;    16'd23346: out <= 16'h0093;    16'd23347: out <= 16'hFC39;
    16'd23348: out <= 16'h0192;    16'd23349: out <= 16'hFE68;    16'd23350: out <= 16'h085D;    16'd23351: out <= 16'h0297;
    16'd23352: out <= 16'h041D;    16'd23353: out <= 16'h000C;    16'd23354: out <= 16'hFF51;    16'd23355: out <= 16'h03A5;
    16'd23356: out <= 16'h0129;    16'd23357: out <= 16'h030D;    16'd23358: out <= 16'hFE24;    16'd23359: out <= 16'hFF4A;
    16'd23360: out <= 16'h0ABD;    16'd23361: out <= 16'hFF2D;    16'd23362: out <= 16'h0A14;    16'd23363: out <= 16'h00B8;
    16'd23364: out <= 16'h03AA;    16'd23365: out <= 16'h0431;    16'd23366: out <= 16'hFD7B;    16'd23367: out <= 16'h0175;
    16'd23368: out <= 16'h0537;    16'd23369: out <= 16'h0AF1;    16'd23370: out <= 16'h07D7;    16'd23371: out <= 16'hFFAE;
    16'd23372: out <= 16'h0492;    16'd23373: out <= 16'h0082;    16'd23374: out <= 16'h0179;    16'd23375: out <= 16'hFD1E;
    16'd23376: out <= 16'h015E;    16'd23377: out <= 16'hFF30;    16'd23378: out <= 16'h02EC;    16'd23379: out <= 16'h0496;
    16'd23380: out <= 16'h0088;    16'd23381: out <= 16'h06B5;    16'd23382: out <= 16'h0964;    16'd23383: out <= 16'hFE30;
    16'd23384: out <= 16'h07E8;    16'd23385: out <= 16'h0A7E;    16'd23386: out <= 16'h00F7;    16'd23387: out <= 16'h04AE;
    16'd23388: out <= 16'h099D;    16'd23389: out <= 16'h0010;    16'd23390: out <= 16'h0068;    16'd23391: out <= 16'h0B63;
    16'd23392: out <= 16'h06A2;    16'd23393: out <= 16'h0799;    16'd23394: out <= 16'h0504;    16'd23395: out <= 16'h0961;
    16'd23396: out <= 16'h0375;    16'd23397: out <= 16'h064A;    16'd23398: out <= 16'hFF7A;    16'd23399: out <= 16'h0847;
    16'd23400: out <= 16'h0401;    16'd23401: out <= 16'h0303;    16'd23402: out <= 16'h014D;    16'd23403: out <= 16'h0525;
    16'd23404: out <= 16'h0A76;    16'd23405: out <= 16'h0479;    16'd23406: out <= 16'h011E;    16'd23407: out <= 16'h097A;
    16'd23408: out <= 16'h03C2;    16'd23409: out <= 16'h063C;    16'd23410: out <= 16'hFC9D;    16'd23411: out <= 16'h05D7;
    16'd23412: out <= 16'h099A;    16'd23413: out <= 16'h0413;    16'd23414: out <= 16'h09F9;    16'd23415: out <= 16'h0486;
    16'd23416: out <= 16'hFFE4;    16'd23417: out <= 16'h04B3;    16'd23418: out <= 16'h01FC;    16'd23419: out <= 16'h012D;
    16'd23420: out <= 16'h0278;    16'd23421: out <= 16'h05B2;    16'd23422: out <= 16'hFF5C;    16'd23423: out <= 16'h0540;
    16'd23424: out <= 16'h03E6;    16'd23425: out <= 16'h093D;    16'd23426: out <= 16'h042D;    16'd23427: out <= 16'h0B6E;
    16'd23428: out <= 16'hFE3A;    16'd23429: out <= 16'h0110;    16'd23430: out <= 16'h08E0;    16'd23431: out <= 16'h0263;
    16'd23432: out <= 16'h065D;    16'd23433: out <= 16'h0649;    16'd23434: out <= 16'h069B;    16'd23435: out <= 16'h08D3;
    16'd23436: out <= 16'hFF8B;    16'd23437: out <= 16'h0394;    16'd23438: out <= 16'h05D2;    16'd23439: out <= 16'h02B4;
    16'd23440: out <= 16'h0012;    16'd23441: out <= 16'hFF59;    16'd23442: out <= 16'hF963;    16'd23443: out <= 16'h0092;
    16'd23444: out <= 16'h03CC;    16'd23445: out <= 16'hFD2D;    16'd23446: out <= 16'hFB9F;    16'd23447: out <= 16'h079F;
    16'd23448: out <= 16'h0082;    16'd23449: out <= 16'h03D2;    16'd23450: out <= 16'h01EE;    16'd23451: out <= 16'hFC15;
    16'd23452: out <= 16'hFF36;    16'd23453: out <= 16'h0039;    16'd23454: out <= 16'h0115;    16'd23455: out <= 16'h011E;
    16'd23456: out <= 16'hFEF5;    16'd23457: out <= 16'h096A;    16'd23458: out <= 16'h06D1;    16'd23459: out <= 16'h0129;
    16'd23460: out <= 16'h0393;    16'd23461: out <= 16'h0C8F;    16'd23462: out <= 16'h01EE;    16'd23463: out <= 16'h093F;
    16'd23464: out <= 16'h008A;    16'd23465: out <= 16'h06FB;    16'd23466: out <= 16'h0D5F;    16'd23467: out <= 16'h0823;
    16'd23468: out <= 16'h0122;    16'd23469: out <= 16'h047E;    16'd23470: out <= 16'h04AD;    16'd23471: out <= 16'h0050;
    16'd23472: out <= 16'h00E8;    16'd23473: out <= 16'h0B95;    16'd23474: out <= 16'h06F5;    16'd23475: out <= 16'hFE69;
    16'd23476: out <= 16'h018F;    16'd23477: out <= 16'h03FD;    16'd23478: out <= 16'h0023;    16'd23479: out <= 16'h023B;
    16'd23480: out <= 16'h05C5;    16'd23481: out <= 16'hFD80;    16'd23482: out <= 16'h06A4;    16'd23483: out <= 16'hF974;
    16'd23484: out <= 16'h0462;    16'd23485: out <= 16'hFADD;    16'd23486: out <= 16'h0576;    16'd23487: out <= 16'h0971;
    16'd23488: out <= 16'h051F;    16'd23489: out <= 16'h05DE;    16'd23490: out <= 16'h0401;    16'd23491: out <= 16'hFCF9;
    16'd23492: out <= 16'h05DC;    16'd23493: out <= 16'h075F;    16'd23494: out <= 16'h03D1;    16'd23495: out <= 16'hFB19;
    16'd23496: out <= 16'h02EC;    16'd23497: out <= 16'h05EB;    16'd23498: out <= 16'hFF05;    16'd23499: out <= 16'h02C7;
    16'd23500: out <= 16'h08EC;    16'd23501: out <= 16'h0704;    16'd23502: out <= 16'h02FD;    16'd23503: out <= 16'h006E;
    16'd23504: out <= 16'h0677;    16'd23505: out <= 16'h03C0;    16'd23506: out <= 16'h01D5;    16'd23507: out <= 16'h078E;
    16'd23508: out <= 16'h03BC;    16'd23509: out <= 16'h05E2;    16'd23510: out <= 16'h03A7;    16'd23511: out <= 16'h047C;
    16'd23512: out <= 16'h02B2;    16'd23513: out <= 16'h074E;    16'd23514: out <= 16'h0843;    16'd23515: out <= 16'h01E2;
    16'd23516: out <= 16'h0237;    16'd23517: out <= 16'h02EE;    16'd23518: out <= 16'h0631;    16'd23519: out <= 16'h0258;
    16'd23520: out <= 16'h04B5;    16'd23521: out <= 16'hFD5E;    16'd23522: out <= 16'h0260;    16'd23523: out <= 16'h00CE;
    16'd23524: out <= 16'h030A;    16'd23525: out <= 16'h0063;    16'd23526: out <= 16'h02B9;    16'd23527: out <= 16'h0114;
    16'd23528: out <= 16'hFF76;    16'd23529: out <= 16'hFFFD;    16'd23530: out <= 16'hFD38;    16'd23531: out <= 16'hFCC8;
    16'd23532: out <= 16'h01E6;    16'd23533: out <= 16'hFE96;    16'd23534: out <= 16'hFB8B;    16'd23535: out <= 16'hFDBE;
    16'd23536: out <= 16'h02BD;    16'd23537: out <= 16'h00E4;    16'd23538: out <= 16'hFBE7;    16'd23539: out <= 16'hFCA2;
    16'd23540: out <= 16'hFB0E;    16'd23541: out <= 16'hFD41;    16'd23542: out <= 16'h04DE;    16'd23543: out <= 16'hFAF9;
    16'd23544: out <= 16'h01DF;    16'd23545: out <= 16'hFE9C;    16'd23546: out <= 16'hFA8D;    16'd23547: out <= 16'hFE9A;
    16'd23548: out <= 16'hFF6E;    16'd23549: out <= 16'h0570;    16'd23550: out <= 16'h006C;    16'd23551: out <= 16'hF89E;
    16'd23552: out <= 16'hFE8E;    16'd23553: out <= 16'h022C;    16'd23554: out <= 16'hFE48;    16'd23555: out <= 16'h0035;
    16'd23556: out <= 16'hFEAD;    16'd23557: out <= 16'h031F;    16'd23558: out <= 16'h01E4;    16'd23559: out <= 16'hFCB2;
    16'd23560: out <= 16'h0168;    16'd23561: out <= 16'h024B;    16'd23562: out <= 16'h0170;    16'd23563: out <= 16'h0631;
    16'd23564: out <= 16'h0252;    16'd23565: out <= 16'hF99E;    16'd23566: out <= 16'hFE87;    16'd23567: out <= 16'h0324;
    16'd23568: out <= 16'h03C0;    16'd23569: out <= 16'h05DE;    16'd23570: out <= 16'hFDCE;    16'd23571: out <= 16'h00D5;
    16'd23572: out <= 16'hFFD6;    16'd23573: out <= 16'hFE3E;    16'd23574: out <= 16'h0129;    16'd23575: out <= 16'h0B2E;
    16'd23576: out <= 16'hFF5E;    16'd23577: out <= 16'hF7E5;    16'd23578: out <= 16'h0130;    16'd23579: out <= 16'hFD91;
    16'd23580: out <= 16'hFFFB;    16'd23581: out <= 16'h01D7;    16'd23582: out <= 16'h0A43;    16'd23583: out <= 16'h01B7;
    16'd23584: out <= 16'h067D;    16'd23585: out <= 16'h0517;    16'd23586: out <= 16'h063D;    16'd23587: out <= 16'h05A7;
    16'd23588: out <= 16'h060F;    16'd23589: out <= 16'h08AA;    16'd23590: out <= 16'h0735;    16'd23591: out <= 16'h0432;
    16'd23592: out <= 16'h001F;    16'd23593: out <= 16'h055B;    16'd23594: out <= 16'hFD3D;    16'd23595: out <= 16'h0533;
    16'd23596: out <= 16'h0D8F;    16'd23597: out <= 16'h03E9;    16'd23598: out <= 16'h0036;    16'd23599: out <= 16'h012B;
    16'd23600: out <= 16'h035B;    16'd23601: out <= 16'h0A65;    16'd23602: out <= 16'h02FE;    16'd23603: out <= 16'h03A0;
    16'd23604: out <= 16'h0536;    16'd23605: out <= 16'hFCB9;    16'd23606: out <= 16'hFED6;    16'd23607: out <= 16'h0F0C;
    16'd23608: out <= 16'h06AF;    16'd23609: out <= 16'h00E7;    16'd23610: out <= 16'h0392;    16'd23611: out <= 16'hFBED;
    16'd23612: out <= 16'h0754;    16'd23613: out <= 16'h0B20;    16'd23614: out <= 16'h041B;    16'd23615: out <= 16'h0158;
    16'd23616: out <= 16'h0596;    16'd23617: out <= 16'h02C0;    16'd23618: out <= 16'h0426;    16'd23619: out <= 16'h0032;
    16'd23620: out <= 16'h06DD;    16'd23621: out <= 16'h058D;    16'd23622: out <= 16'h03FF;    16'd23623: out <= 16'hFE64;
    16'd23624: out <= 16'h03A7;    16'd23625: out <= 16'h0520;    16'd23626: out <= 16'h02E2;    16'd23627: out <= 16'h0887;
    16'd23628: out <= 16'h0399;    16'd23629: out <= 16'h0256;    16'd23630: out <= 16'h0D5C;    16'd23631: out <= 16'hFCFE;
    16'd23632: out <= 16'hFF36;    16'd23633: out <= 16'h03E0;    16'd23634: out <= 16'h047A;    16'd23635: out <= 16'h0422;
    16'd23636: out <= 16'h010D;    16'd23637: out <= 16'hFEDB;    16'd23638: out <= 16'h0C35;    16'd23639: out <= 16'h017B;
    16'd23640: out <= 16'h0A8B;    16'd23641: out <= 16'h0435;    16'd23642: out <= 16'hFDF1;    16'd23643: out <= 16'h00EC;
    16'd23644: out <= 16'h04C7;    16'd23645: out <= 16'h085C;    16'd23646: out <= 16'hFFBB;    16'd23647: out <= 16'hFC12;
    16'd23648: out <= 16'h0420;    16'd23649: out <= 16'hFEB2;    16'd23650: out <= 16'h0C09;    16'd23651: out <= 16'h0330;
    16'd23652: out <= 16'h03EC;    16'd23653: out <= 16'h07F7;    16'd23654: out <= 16'h02CF;    16'd23655: out <= 16'hFDCD;
    16'd23656: out <= 16'h0172;    16'd23657: out <= 16'h0055;    16'd23658: out <= 16'h050B;    16'd23659: out <= 16'h08DF;
    16'd23660: out <= 16'h0852;    16'd23661: out <= 16'h02D6;    16'd23662: out <= 16'h0526;    16'd23663: out <= 16'h0377;
    16'd23664: out <= 16'hFFCF;    16'd23665: out <= 16'h0415;    16'd23666: out <= 16'h0543;    16'd23667: out <= 16'h0385;
    16'd23668: out <= 16'h0481;    16'd23669: out <= 16'h07B6;    16'd23670: out <= 16'hFF26;    16'd23671: out <= 16'h0379;
    16'd23672: out <= 16'h00BE;    16'd23673: out <= 16'h0737;    16'd23674: out <= 16'h0840;    16'd23675: out <= 16'hFEAE;
    16'd23676: out <= 16'h00FE;    16'd23677: out <= 16'h071B;    16'd23678: out <= 16'h092B;    16'd23679: out <= 16'hFAE3;
    16'd23680: out <= 16'h04D3;    16'd23681: out <= 16'h0115;    16'd23682: out <= 16'hFE3E;    16'd23683: out <= 16'h0544;
    16'd23684: out <= 16'h0150;    16'd23685: out <= 16'h0268;    16'd23686: out <= 16'h076F;    16'd23687: out <= 16'hFECC;
    16'd23688: out <= 16'h0354;    16'd23689: out <= 16'h008A;    16'd23690: out <= 16'h0426;    16'd23691: out <= 16'hFF64;
    16'd23692: out <= 16'h05EE;    16'd23693: out <= 16'h045C;    16'd23694: out <= 16'h0442;    16'd23695: out <= 16'h02E0;
    16'd23696: out <= 16'hF6B6;    16'd23697: out <= 16'h0192;    16'd23698: out <= 16'h00AD;    16'd23699: out <= 16'h00F6;
    16'd23700: out <= 16'hFE58;    16'd23701: out <= 16'h01A6;    16'd23702: out <= 16'hFD18;    16'd23703: out <= 16'hFCED;
    16'd23704: out <= 16'h0244;    16'd23705: out <= 16'h022E;    16'd23706: out <= 16'h0519;    16'd23707: out <= 16'h02F9;
    16'd23708: out <= 16'h06F9;    16'd23709: out <= 16'hFA9C;    16'd23710: out <= 16'h06AC;    16'd23711: out <= 16'h0036;
    16'd23712: out <= 16'hFE36;    16'd23713: out <= 16'h0606;    16'd23714: out <= 16'h0180;    16'd23715: out <= 16'hFCE4;
    16'd23716: out <= 16'h0C0D;    16'd23717: out <= 16'h06FE;    16'd23718: out <= 16'h04DE;    16'd23719: out <= 16'h0502;
    16'd23720: out <= 16'h03BC;    16'd23721: out <= 16'h0936;    16'd23722: out <= 16'h000E;    16'd23723: out <= 16'h04EF;
    16'd23724: out <= 16'h0254;    16'd23725: out <= 16'h076F;    16'd23726: out <= 16'h00F4;    16'd23727: out <= 16'h05EA;
    16'd23728: out <= 16'hFF82;    16'd23729: out <= 16'h02F2;    16'd23730: out <= 16'h05FA;    16'd23731: out <= 16'h050B;
    16'd23732: out <= 16'h08B1;    16'd23733: out <= 16'h0D3D;    16'd23734: out <= 16'h0AE4;    16'd23735: out <= 16'h0654;
    16'd23736: out <= 16'h03AD;    16'd23737: out <= 16'h06A4;    16'd23738: out <= 16'hFE54;    16'd23739: out <= 16'h04D9;
    16'd23740: out <= 16'h06C3;    16'd23741: out <= 16'h0439;    16'd23742: out <= 16'h082E;    16'd23743: out <= 16'h0051;
    16'd23744: out <= 16'h0782;    16'd23745: out <= 16'h045B;    16'd23746: out <= 16'h0434;    16'd23747: out <= 16'h0636;
    16'd23748: out <= 16'h0882;    16'd23749: out <= 16'h0482;    16'd23750: out <= 16'h02C2;    16'd23751: out <= 16'h030F;
    16'd23752: out <= 16'h02C0;    16'd23753: out <= 16'hFD45;    16'd23754: out <= 16'h02B6;    16'd23755: out <= 16'h060D;
    16'd23756: out <= 16'hFF2A;    16'd23757: out <= 16'h09D2;    16'd23758: out <= 16'h00DD;    16'd23759: out <= 16'h0144;
    16'd23760: out <= 16'h0493;    16'd23761: out <= 16'h02FD;    16'd23762: out <= 16'h047D;    16'd23763: out <= 16'h0223;
    16'd23764: out <= 16'h044F;    16'd23765: out <= 16'h0492;    16'd23766: out <= 16'h019F;    16'd23767: out <= 16'h0002;
    16'd23768: out <= 16'h042B;    16'd23769: out <= 16'h039E;    16'd23770: out <= 16'h0942;    16'd23771: out <= 16'hFEF1;
    16'd23772: out <= 16'h03E1;    16'd23773: out <= 16'hFE59;    16'd23774: out <= 16'hF97B;    16'd23775: out <= 16'h07AF;
    16'd23776: out <= 16'hF9EC;    16'd23777: out <= 16'hF908;    16'd23778: out <= 16'h0740;    16'd23779: out <= 16'h0121;
    16'd23780: out <= 16'hFC36;    16'd23781: out <= 16'hF646;    16'd23782: out <= 16'h0014;    16'd23783: out <= 16'h0292;
    16'd23784: out <= 16'hFA85;    16'd23785: out <= 16'h040B;    16'd23786: out <= 16'h01F2;    16'd23787: out <= 16'h01BC;
    16'd23788: out <= 16'hFF9F;    16'd23789: out <= 16'hFE48;    16'd23790: out <= 16'hFDA6;    16'd23791: out <= 16'hFE1B;
    16'd23792: out <= 16'hFE78;    16'd23793: out <= 16'h03EB;    16'd23794: out <= 16'hFDC5;    16'd23795: out <= 16'h0220;
    16'd23796: out <= 16'hFF15;    16'd23797: out <= 16'hFAF4;    16'd23798: out <= 16'h038F;    16'd23799: out <= 16'hFCF5;
    16'd23800: out <= 16'hFBA2;    16'd23801: out <= 16'h0612;    16'd23802: out <= 16'hFD52;    16'd23803: out <= 16'h0763;
    16'd23804: out <= 16'hFF37;    16'd23805: out <= 16'h0416;    16'd23806: out <= 16'hFF0B;    16'd23807: out <= 16'hFEFD;
    16'd23808: out <= 16'h0121;    16'd23809: out <= 16'hF7E4;    16'd23810: out <= 16'h05B3;    16'd23811: out <= 16'hFB6B;
    16'd23812: out <= 16'hFDE1;    16'd23813: out <= 16'h0407;    16'd23814: out <= 16'hFFDD;    16'd23815: out <= 16'h0574;
    16'd23816: out <= 16'hFF51;    16'd23817: out <= 16'hFC2A;    16'd23818: out <= 16'h023F;    16'd23819: out <= 16'h0362;
    16'd23820: out <= 16'hFA77;    16'd23821: out <= 16'hFF3E;    16'd23822: out <= 16'hFCB4;    16'd23823: out <= 16'h032A;
    16'd23824: out <= 16'h056A;    16'd23825: out <= 16'h040B;    16'd23826: out <= 16'hFA7B;    16'd23827: out <= 16'h00F5;
    16'd23828: out <= 16'h0332;    16'd23829: out <= 16'hFB22;    16'd23830: out <= 16'hFE11;    16'd23831: out <= 16'h0391;
    16'd23832: out <= 16'h05F1;    16'd23833: out <= 16'h0377;    16'd23834: out <= 16'hFA13;    16'd23835: out <= 16'hFAEE;
    16'd23836: out <= 16'h00F2;    16'd23837: out <= 16'h0AB3;    16'd23838: out <= 16'hFC66;    16'd23839: out <= 16'h00E0;
    16'd23840: out <= 16'h062E;    16'd23841: out <= 16'h028C;    16'd23842: out <= 16'h0BB7;    16'd23843: out <= 16'hFF8C;
    16'd23844: out <= 16'h0167;    16'd23845: out <= 16'h042E;    16'd23846: out <= 16'hFD33;    16'd23847: out <= 16'h03C0;
    16'd23848: out <= 16'h01DE;    16'd23849: out <= 16'h0AC1;    16'd23850: out <= 16'h0337;    16'd23851: out <= 16'h0094;
    16'd23852: out <= 16'h0779;    16'd23853: out <= 16'h010D;    16'd23854: out <= 16'h0142;    16'd23855: out <= 16'hFE1A;
    16'd23856: out <= 16'h0BC7;    16'd23857: out <= 16'h0136;    16'd23858: out <= 16'h0961;    16'd23859: out <= 16'h03B3;
    16'd23860: out <= 16'h05D7;    16'd23861: out <= 16'h02CF;    16'd23862: out <= 16'h02E7;    16'd23863: out <= 16'h03B4;
    16'd23864: out <= 16'hFE67;    16'd23865: out <= 16'h03DF;    16'd23866: out <= 16'h036D;    16'd23867: out <= 16'h028E;
    16'd23868: out <= 16'h063A;    16'd23869: out <= 16'h062B;    16'd23870: out <= 16'h0009;    16'd23871: out <= 16'h08BD;
    16'd23872: out <= 16'h04CF;    16'd23873: out <= 16'h0742;    16'd23874: out <= 16'hFCCF;    16'd23875: out <= 16'hFF36;
    16'd23876: out <= 16'h0516;    16'd23877: out <= 16'h04C0;    16'd23878: out <= 16'hFC89;    16'd23879: out <= 16'h0BBF;
    16'd23880: out <= 16'h03D9;    16'd23881: out <= 16'h0040;    16'd23882: out <= 16'h00F0;    16'd23883: out <= 16'h08CA;
    16'd23884: out <= 16'h018D;    16'd23885: out <= 16'h0257;    16'd23886: out <= 16'h0A16;    16'd23887: out <= 16'h01C1;
    16'd23888: out <= 16'h039A;    16'd23889: out <= 16'h0288;    16'd23890: out <= 16'h005E;    16'd23891: out <= 16'h04D6;
    16'd23892: out <= 16'hFEB3;    16'd23893: out <= 16'h04AD;    16'd23894: out <= 16'h059D;    16'd23895: out <= 16'h073A;
    16'd23896: out <= 16'h058F;    16'd23897: out <= 16'h0133;    16'd23898: out <= 16'h02F7;    16'd23899: out <= 16'hFEFB;
    16'd23900: out <= 16'h0380;    16'd23901: out <= 16'h04EF;    16'd23902: out <= 16'h04DE;    16'd23903: out <= 16'h09EF;
    16'd23904: out <= 16'hFF5D;    16'd23905: out <= 16'h060A;    16'd23906: out <= 16'h0B4F;    16'd23907: out <= 16'h036C;
    16'd23908: out <= 16'h04C1;    16'd23909: out <= 16'h0651;    16'd23910: out <= 16'hFBB2;    16'd23911: out <= 16'h0106;
    16'd23912: out <= 16'h084C;    16'd23913: out <= 16'h0900;    16'd23914: out <= 16'h01AC;    16'd23915: out <= 16'h027F;
    16'd23916: out <= 16'h0A63;    16'd23917: out <= 16'h04BF;    16'd23918: out <= 16'h033B;    16'd23919: out <= 16'h05E7;
    16'd23920: out <= 16'h099F;    16'd23921: out <= 16'h0616;    16'd23922: out <= 16'hFF35;    16'd23923: out <= 16'h026E;
    16'd23924: out <= 16'h0373;    16'd23925: out <= 16'h0569;    16'd23926: out <= 16'hFFED;    16'd23927: out <= 16'hFED8;
    16'd23928: out <= 16'h047F;    16'd23929: out <= 16'h00BF;    16'd23930: out <= 16'hFF4C;    16'd23931: out <= 16'hFDEE;
    16'd23932: out <= 16'hFF56;    16'd23933: out <= 16'h0D04;    16'd23934: out <= 16'h02F1;    16'd23935: out <= 16'h031F;
    16'd23936: out <= 16'h04F2;    16'd23937: out <= 16'h02F2;    16'd23938: out <= 16'h067F;    16'd23939: out <= 16'h049F;
    16'd23940: out <= 16'h06D1;    16'd23941: out <= 16'h0A0A;    16'd23942: out <= 16'h0306;    16'd23943: out <= 16'h0686;
    16'd23944: out <= 16'hFF0E;    16'd23945: out <= 16'h075D;    16'd23946: out <= 16'h0173;    16'd23947: out <= 16'h0518;
    16'd23948: out <= 16'h001C;    16'd23949: out <= 16'h0403;    16'd23950: out <= 16'h0894;    16'd23951: out <= 16'hF92F;
    16'd23952: out <= 16'h0068;    16'd23953: out <= 16'h03FB;    16'd23954: out <= 16'h06D3;    16'd23955: out <= 16'hFE8B;
    16'd23956: out <= 16'h08F1;    16'd23957: out <= 16'h02AE;    16'd23958: out <= 16'h076A;    16'd23959: out <= 16'hFF66;
    16'd23960: out <= 16'hFED3;    16'd23961: out <= 16'hFA58;    16'd23962: out <= 16'hFB7F;    16'd23963: out <= 16'h019E;
    16'd23964: out <= 16'hF9E1;    16'd23965: out <= 16'h0370;    16'd23966: out <= 16'hFD43;    16'd23967: out <= 16'hFFEF;
    16'd23968: out <= 16'h0237;    16'd23969: out <= 16'h053D;    16'd23970: out <= 16'h08AD;    16'd23971: out <= 16'h0311;
    16'd23972: out <= 16'h00E8;    16'd23973: out <= 16'h08BB;    16'd23974: out <= 16'h06C9;    16'd23975: out <= 16'hFDE7;
    16'd23976: out <= 16'hFE29;    16'd23977: out <= 16'h011C;    16'd23978: out <= 16'h0216;    16'd23979: out <= 16'h0535;
    16'd23980: out <= 16'h03D2;    16'd23981: out <= 16'h03DB;    16'd23982: out <= 16'h0566;    16'd23983: out <= 16'h0145;
    16'd23984: out <= 16'h03AF;    16'd23985: out <= 16'h0874;    16'd23986: out <= 16'h033E;    16'd23987: out <= 16'h025A;
    16'd23988: out <= 16'h0068;    16'd23989: out <= 16'h0416;    16'd23990: out <= 16'h0730;    16'd23991: out <= 16'h09CB;
    16'd23992: out <= 16'hFD18;    16'd23993: out <= 16'h00B3;    16'd23994: out <= 16'h03E5;    16'd23995: out <= 16'h05AE;
    16'd23996: out <= 16'h06C4;    16'd23997: out <= 16'hFB87;    16'd23998: out <= 16'h0301;    16'd23999: out <= 16'h0273;
    16'd24000: out <= 16'h0094;    16'd24001: out <= 16'hFF05;    16'd24002: out <= 16'h0109;    16'd24003: out <= 16'h0378;
    16'd24004: out <= 16'h087C;    16'd24005: out <= 16'h052A;    16'd24006: out <= 16'h01EC;    16'd24007: out <= 16'h04D1;
    16'd24008: out <= 16'h0478;    16'd24009: out <= 16'h07AF;    16'd24010: out <= 16'h0470;    16'd24011: out <= 16'h0699;
    16'd24012: out <= 16'h05F4;    16'd24013: out <= 16'h036E;    16'd24014: out <= 16'h00E6;    16'd24015: out <= 16'h0566;
    16'd24016: out <= 16'h018E;    16'd24017: out <= 16'h01B0;    16'd24018: out <= 16'h0246;    16'd24019: out <= 16'h07A5;
    16'd24020: out <= 16'hFFC6;    16'd24021: out <= 16'h05B3;    16'd24022: out <= 16'h008E;    16'd24023: out <= 16'h047B;
    16'd24024: out <= 16'h09A2;    16'd24025: out <= 16'hFE4E;    16'd24026: out <= 16'hFF53;    16'd24027: out <= 16'h0156;
    16'd24028: out <= 16'hFC78;    16'd24029: out <= 16'h0691;    16'd24030: out <= 16'h00AD;    16'd24031: out <= 16'hFF8D;
    16'd24032: out <= 16'hFD9B;    16'd24033: out <= 16'hFB66;    16'd24034: out <= 16'h01C2;    16'd24035: out <= 16'h0447;
    16'd24036: out <= 16'hFD3C;    16'd24037: out <= 16'h0029;    16'd24038: out <= 16'h0457;    16'd24039: out <= 16'h02D9;
    16'd24040: out <= 16'hFE38;    16'd24041: out <= 16'h0088;    16'd24042: out <= 16'h0053;    16'd24043: out <= 16'hFB3F;
    16'd24044: out <= 16'hF79B;    16'd24045: out <= 16'hFF69;    16'd24046: out <= 16'hF9E7;    16'd24047: out <= 16'h040A;
    16'd24048: out <= 16'hFFB4;    16'd24049: out <= 16'hFE06;    16'd24050: out <= 16'hFCAC;    16'd24051: out <= 16'h00C6;
    16'd24052: out <= 16'h055A;    16'd24053: out <= 16'hF846;    16'd24054: out <= 16'hF8A8;    16'd24055: out <= 16'hFC95;
    16'd24056: out <= 16'h0010;    16'd24057: out <= 16'hFA64;    16'd24058: out <= 16'h03A7;    16'd24059: out <= 16'hFBFE;
    16'd24060: out <= 16'hFE30;    16'd24061: out <= 16'h10F8;    16'd24062: out <= 16'h0591;    16'd24063: out <= 16'h0084;
    16'd24064: out <= 16'hFD49;    16'd24065: out <= 16'hFCEA;    16'd24066: out <= 16'h0000;    16'd24067: out <= 16'hFED8;
    16'd24068: out <= 16'hFDEE;    16'd24069: out <= 16'h0693;    16'd24070: out <= 16'h04E9;    16'd24071: out <= 16'h02B9;
    16'd24072: out <= 16'hFE44;    16'd24073: out <= 16'h031D;    16'd24074: out <= 16'h063D;    16'd24075: out <= 16'h0085;
    16'd24076: out <= 16'hFF33;    16'd24077: out <= 16'h0396;    16'd24078: out <= 16'h02FC;    16'd24079: out <= 16'h062E;
    16'd24080: out <= 16'hFE83;    16'd24081: out <= 16'hFB90;    16'd24082: out <= 16'hFE4B;    16'd24083: out <= 16'hFDDC;
    16'd24084: out <= 16'hFF6A;    16'd24085: out <= 16'h02C0;    16'd24086: out <= 16'hFFCB;    16'd24087: out <= 16'h02B4;
    16'd24088: out <= 16'hFFC5;    16'd24089: out <= 16'h0565;    16'd24090: out <= 16'h000F;    16'd24091: out <= 16'h0136;
    16'd24092: out <= 16'h0307;    16'd24093: out <= 16'h0425;    16'd24094: out <= 16'h04B7;    16'd24095: out <= 16'h0410;
    16'd24096: out <= 16'hFE4F;    16'd24097: out <= 16'h04D2;    16'd24098: out <= 16'h023C;    16'd24099: out <= 16'h0252;
    16'd24100: out <= 16'h06CC;    16'd24101: out <= 16'h04A6;    16'd24102: out <= 16'h0459;    16'd24103: out <= 16'h03B2;
    16'd24104: out <= 16'h0C18;    16'd24105: out <= 16'h003D;    16'd24106: out <= 16'h0845;    16'd24107: out <= 16'h04A2;
    16'd24108: out <= 16'h0A2E;    16'd24109: out <= 16'h0359;    16'd24110: out <= 16'h0863;    16'd24111: out <= 16'h0022;
    16'd24112: out <= 16'h0A51;    16'd24113: out <= 16'h054F;    16'd24114: out <= 16'h03FF;    16'd24115: out <= 16'h0671;
    16'd24116: out <= 16'h09C5;    16'd24117: out <= 16'h01E9;    16'd24118: out <= 16'hFF48;    16'd24119: out <= 16'h017B;
    16'd24120: out <= 16'h04C8;    16'd24121: out <= 16'hFF7C;    16'd24122: out <= 16'h057A;    16'd24123: out <= 16'h031B;
    16'd24124: out <= 16'h0191;    16'd24125: out <= 16'h0769;    16'd24126: out <= 16'h0936;    16'd24127: out <= 16'h06FB;
    16'd24128: out <= 16'hFFED;    16'd24129: out <= 16'h013F;    16'd24130: out <= 16'h0D6C;    16'd24131: out <= 16'h0518;
    16'd24132: out <= 16'h0045;    16'd24133: out <= 16'h0597;    16'd24134: out <= 16'h09A3;    16'd24135: out <= 16'h02C7;
    16'd24136: out <= 16'h09D0;    16'd24137: out <= 16'h035D;    16'd24138: out <= 16'h063C;    16'd24139: out <= 16'h0744;
    16'd24140: out <= 16'h02CF;    16'd24141: out <= 16'h0714;    16'd24142: out <= 16'h0086;    16'd24143: out <= 16'h003A;
    16'd24144: out <= 16'hFC6D;    16'd24145: out <= 16'hFB8E;    16'd24146: out <= 16'h0346;    16'd24147: out <= 16'h0452;
    16'd24148: out <= 16'hFF47;    16'd24149: out <= 16'h0268;    16'd24150: out <= 16'h05C4;    16'd24151: out <= 16'h067F;
    16'd24152: out <= 16'h024F;    16'd24153: out <= 16'h0AE9;    16'd24154: out <= 16'h06A9;    16'd24155: out <= 16'h098A;
    16'd24156: out <= 16'hFA93;    16'd24157: out <= 16'h00C7;    16'd24158: out <= 16'h0590;    16'd24159: out <= 16'hFB5B;
    16'd24160: out <= 16'h00B3;    16'd24161: out <= 16'h033B;    16'd24162: out <= 16'h0389;    16'd24163: out <= 16'h0100;
    16'd24164: out <= 16'h0278;    16'd24165: out <= 16'h0718;    16'd24166: out <= 16'h0933;    16'd24167: out <= 16'h096C;
    16'd24168: out <= 16'h033F;    16'd24169: out <= 16'h0208;    16'd24170: out <= 16'h030F;    16'd24171: out <= 16'h082A;
    16'd24172: out <= 16'h06D5;    16'd24173: out <= 16'h0314;    16'd24174: out <= 16'h0262;    16'd24175: out <= 16'h0484;
    16'd24176: out <= 16'h0135;    16'd24177: out <= 16'h03BC;    16'd24178: out <= 16'h0B7F;    16'd24179: out <= 16'h04DF;
    16'd24180: out <= 16'h00A5;    16'd24181: out <= 16'h02AD;    16'd24182: out <= 16'h023B;    16'd24183: out <= 16'h0260;
    16'd24184: out <= 16'h0789;    16'd24185: out <= 16'h087F;    16'd24186: out <= 16'h0779;    16'd24187: out <= 16'h0C22;
    16'd24188: out <= 16'h0521;    16'd24189: out <= 16'h089B;    16'd24190: out <= 16'h0656;    16'd24191: out <= 16'h061A;
    16'd24192: out <= 16'h060B;    16'd24193: out <= 16'h0724;    16'd24194: out <= 16'h04F5;    16'd24195: out <= 16'h0155;
    16'd24196: out <= 16'h02B4;    16'd24197: out <= 16'h00FF;    16'd24198: out <= 16'h07B9;    16'd24199: out <= 16'hFCA1;
    16'd24200: out <= 16'h08E7;    16'd24201: out <= 16'h040C;    16'd24202: out <= 16'h0404;    16'd24203: out <= 16'h03D4;
    16'd24204: out <= 16'h0CED;    16'd24205: out <= 16'hFF37;    16'd24206: out <= 16'hF9C4;    16'd24207: out <= 16'h038C;
    16'd24208: out <= 16'hFFD1;    16'd24209: out <= 16'h0099;    16'd24210: out <= 16'hFA50;    16'd24211: out <= 16'hFEDE;
    16'd24212: out <= 16'hFBBF;    16'd24213: out <= 16'hF8F7;    16'd24214: out <= 16'h0439;    16'd24215: out <= 16'hFF90;
    16'd24216: out <= 16'h04D3;    16'd24217: out <= 16'h0268;    16'd24218: out <= 16'hFE54;    16'd24219: out <= 16'h0421;
    16'd24220: out <= 16'hFF87;    16'd24221: out <= 16'hFFE0;    16'd24222: out <= 16'h0155;    16'd24223: out <= 16'h0857;
    16'd24224: out <= 16'hFE2D;    16'd24225: out <= 16'hFEC3;    16'd24226: out <= 16'h02F6;    16'd24227: out <= 16'h05D0;
    16'd24228: out <= 16'h0698;    16'd24229: out <= 16'h02BB;    16'd24230: out <= 16'h080C;    16'd24231: out <= 16'h06F2;
    16'd24232: out <= 16'h05B2;    16'd24233: out <= 16'h0982;    16'd24234: out <= 16'h0627;    16'd24235: out <= 16'h025B;
    16'd24236: out <= 16'h0826;    16'd24237: out <= 16'h0204;    16'd24238: out <= 16'h06AE;    16'd24239: out <= 16'hFFAD;
    16'd24240: out <= 16'h0E85;    16'd24241: out <= 16'h08BC;    16'd24242: out <= 16'h03B2;    16'd24243: out <= 16'h0CF9;
    16'd24244: out <= 16'h022A;    16'd24245: out <= 16'h017D;    16'd24246: out <= 16'h0450;    16'd24247: out <= 16'h096A;
    16'd24248: out <= 16'h0C14;    16'd24249: out <= 16'hFEB4;    16'd24250: out <= 16'h06EF;    16'd24251: out <= 16'h02B3;
    16'd24252: out <= 16'h08F4;    16'd24253: out <= 16'h0A5B;    16'd24254: out <= 16'h0706;    16'd24255: out <= 16'h04A0;
    16'd24256: out <= 16'h08F5;    16'd24257: out <= 16'hF89B;    16'd24258: out <= 16'hFC48;    16'd24259: out <= 16'h0017;
    16'd24260: out <= 16'h0485;    16'd24261: out <= 16'h0499;    16'd24262: out <= 16'hFBE2;    16'd24263: out <= 16'h0745;
    16'd24264: out <= 16'h00B7;    16'd24265: out <= 16'h0820;    16'd24266: out <= 16'h095A;    16'd24267: out <= 16'h00E2;
    16'd24268: out <= 16'h07F4;    16'd24269: out <= 16'h0B06;    16'd24270: out <= 16'h0600;    16'd24271: out <= 16'h03EC;
    16'd24272: out <= 16'h0245;    16'd24273: out <= 16'h02B3;    16'd24274: out <= 16'h041D;    16'd24275: out <= 16'hFF90;
    16'd24276: out <= 16'h0720;    16'd24277: out <= 16'h057E;    16'd24278: out <= 16'hFC9A;    16'd24279: out <= 16'h03EE;
    16'd24280: out <= 16'hFD9C;    16'd24281: out <= 16'h03A6;    16'd24282: out <= 16'h03C7;    16'd24283: out <= 16'h02C2;
    16'd24284: out <= 16'h08EE;    16'd24285: out <= 16'h01F5;    16'd24286: out <= 16'h0358;    16'd24287: out <= 16'hFEC4;
    16'd24288: out <= 16'hFEBA;    16'd24289: out <= 16'hFF73;    16'd24290: out <= 16'h008E;    16'd24291: out <= 16'hFCCF;
    16'd24292: out <= 16'hFFEA;    16'd24293: out <= 16'hFD9A;    16'd24294: out <= 16'h03A0;    16'd24295: out <= 16'h0015;
    16'd24296: out <= 16'h00FE;    16'd24297: out <= 16'hFE2D;    16'd24298: out <= 16'h00F5;    16'd24299: out <= 16'h026E;
    16'd24300: out <= 16'h0147;    16'd24301: out <= 16'h012F;    16'd24302: out <= 16'h05B0;    16'd24303: out <= 16'h02F6;
    16'd24304: out <= 16'h0852;    16'd24305: out <= 16'h020C;    16'd24306: out <= 16'hFF4D;    16'd24307: out <= 16'h001F;
    16'd24308: out <= 16'hFAEF;    16'd24309: out <= 16'h001B;    16'd24310: out <= 16'h004A;    16'd24311: out <= 16'hFF47;
    16'd24312: out <= 16'hFAD9;    16'd24313: out <= 16'h00AE;    16'd24314: out <= 16'hF93B;    16'd24315: out <= 16'hFFD6;
    16'd24316: out <= 16'h045C;    16'd24317: out <= 16'h00E2;    16'd24318: out <= 16'h0698;    16'd24319: out <= 16'h0355;
    16'd24320: out <= 16'h029B;    16'd24321: out <= 16'h021D;    16'd24322: out <= 16'h02D5;    16'd24323: out <= 16'hFF55;
    16'd24324: out <= 16'h0119;    16'd24325: out <= 16'h01E8;    16'd24326: out <= 16'h069F;    16'd24327: out <= 16'h0049;
    16'd24328: out <= 16'h039F;    16'd24329: out <= 16'h05CB;    16'd24330: out <= 16'hFD5D;    16'd24331: out <= 16'hFB48;
    16'd24332: out <= 16'hFAF5;    16'd24333: out <= 16'hFD46;    16'd24334: out <= 16'hFC0C;    16'd24335: out <= 16'hFCC1;
    16'd24336: out <= 16'h0225;    16'd24337: out <= 16'hF97D;    16'd24338: out <= 16'h0835;    16'd24339: out <= 16'hFDD9;
    16'd24340: out <= 16'hFEDA;    16'd24341: out <= 16'hFFDA;    16'd24342: out <= 16'h0A4D;    16'd24343: out <= 16'hF8D7;
    16'd24344: out <= 16'hFF56;    16'd24345: out <= 16'h0187;    16'd24346: out <= 16'hFDB2;    16'd24347: out <= 16'h013C;
    16'd24348: out <= 16'h02F8;    16'd24349: out <= 16'h0340;    16'd24350: out <= 16'h0471;    16'd24351: out <= 16'h03D0;
    16'd24352: out <= 16'h052F;    16'd24353: out <= 16'h0342;    16'd24354: out <= 16'h0669;    16'd24355: out <= 16'h02D0;
    16'd24356: out <= 16'h01A9;    16'd24357: out <= 16'hFDEE;    16'd24358: out <= 16'h06FA;    16'd24359: out <= 16'hFD94;
    16'd24360: out <= 16'h087A;    16'd24361: out <= 16'h05B8;    16'd24362: out <= 16'hFD46;    16'd24363: out <= 16'h0280;
    16'd24364: out <= 16'h03C9;    16'd24365: out <= 16'hFFE3;    16'd24366: out <= 16'h04DA;    16'd24367: out <= 16'hFF15;
    16'd24368: out <= 16'h0435;    16'd24369: out <= 16'h0430;    16'd24370: out <= 16'h084E;    16'd24371: out <= 16'h0CEF;
    16'd24372: out <= 16'h0367;    16'd24373: out <= 16'h0406;    16'd24374: out <= 16'hFEE8;    16'd24375: out <= 16'hFF1C;
    16'd24376: out <= 16'hFF66;    16'd24377: out <= 16'hFCBB;    16'd24378: out <= 16'hFDC0;    16'd24379: out <= 16'h03DC;
    16'd24380: out <= 16'hFD56;    16'd24381: out <= 16'h0664;    16'd24382: out <= 16'h0459;    16'd24383: out <= 16'hFF45;
    16'd24384: out <= 16'h0003;    16'd24385: out <= 16'h0468;    16'd24386: out <= 16'h03ED;    16'd24387: out <= 16'h05FB;
    16'd24388: out <= 16'h01B6;    16'd24389: out <= 16'h03F0;    16'd24390: out <= 16'h04AF;    16'd24391: out <= 16'h018D;
    16'd24392: out <= 16'h084A;    16'd24393: out <= 16'h0220;    16'd24394: out <= 16'hFF42;    16'd24395: out <= 16'hFF19;
    16'd24396: out <= 16'h0432;    16'd24397: out <= 16'hFA5A;    16'd24398: out <= 16'h04EC;    16'd24399: out <= 16'h0895;
    16'd24400: out <= 16'h0727;    16'd24401: out <= 16'h04EE;    16'd24402: out <= 16'hFD32;    16'd24403: out <= 16'h0504;
    16'd24404: out <= 16'h049D;    16'd24405: out <= 16'h0812;    16'd24406: out <= 16'h0813;    16'd24407: out <= 16'h02B8;
    16'd24408: out <= 16'h091D;    16'd24409: out <= 16'h0693;    16'd24410: out <= 16'hFF5C;    16'd24411: out <= 16'hFEA5;
    16'd24412: out <= 16'hFFAE;    16'd24413: out <= 16'hF880;    16'd24414: out <= 16'h05DC;    16'd24415: out <= 16'h00F9;
    16'd24416: out <= 16'hFE6E;    16'd24417: out <= 16'hFAEA;    16'd24418: out <= 16'hFE5B;    16'd24419: out <= 16'hFD3A;
    16'd24420: out <= 16'hFDC2;    16'd24421: out <= 16'h0815;    16'd24422: out <= 16'h08CE;    16'd24423: out <= 16'h05E5;
    16'd24424: out <= 16'h06A9;    16'd24425: out <= 16'h03BC;    16'd24426: out <= 16'h0543;    16'd24427: out <= 16'h0544;
    16'd24428: out <= 16'h098D;    16'd24429: out <= 16'hFF39;    16'd24430: out <= 16'h064E;    16'd24431: out <= 16'h0404;
    16'd24432: out <= 16'h08B1;    16'd24433: out <= 16'hFCF9;    16'd24434: out <= 16'h022E;    16'd24435: out <= 16'h02A2;
    16'd24436: out <= 16'hFD62;    16'd24437: out <= 16'hFFA0;    16'd24438: out <= 16'h0774;    16'd24439: out <= 16'h02C2;
    16'd24440: out <= 16'h06CD;    16'd24441: out <= 16'h00F8;    16'd24442: out <= 16'h01BF;    16'd24443: out <= 16'h0728;
    16'd24444: out <= 16'h05F6;    16'd24445: out <= 16'hFEF8;    16'd24446: out <= 16'hFCFE;    16'd24447: out <= 16'hFFF2;
    16'd24448: out <= 16'h0072;    16'd24449: out <= 16'h000A;    16'd24450: out <= 16'h04C0;    16'd24451: out <= 16'h00CA;
    16'd24452: out <= 16'h0781;    16'd24453: out <= 16'h0365;    16'd24454: out <= 16'hFDF2;    16'd24455: out <= 16'h044B;
    16'd24456: out <= 16'h0B1F;    16'd24457: out <= 16'h0449;    16'd24458: out <= 16'hFC3C;    16'd24459: out <= 16'h053F;
    16'd24460: out <= 16'h0081;    16'd24461: out <= 16'hF8FD;    16'd24462: out <= 16'hFC74;    16'd24463: out <= 16'h00BA;
    16'd24464: out <= 16'hFD02;    16'd24465: out <= 16'h013D;    16'd24466: out <= 16'h031A;    16'd24467: out <= 16'hFF0B;
    16'd24468: out <= 16'h03E1;    16'd24469: out <= 16'h0003;    16'd24470: out <= 16'h044A;    16'd24471: out <= 16'hFBED;
    16'd24472: out <= 16'hFCDA;    16'd24473: out <= 16'hFF43;    16'd24474: out <= 16'hFE08;    16'd24475: out <= 16'hFA0E;
    16'd24476: out <= 16'h046F;    16'd24477: out <= 16'h0887;    16'd24478: out <= 16'hFB51;    16'd24479: out <= 16'h0512;
    16'd24480: out <= 16'h081D;    16'd24481: out <= 16'h01F7;    16'd24482: out <= 16'h03AA;    16'd24483: out <= 16'hFF33;
    16'd24484: out <= 16'h09CD;    16'd24485: out <= 16'h0131;    16'd24486: out <= 16'h00A9;    16'd24487: out <= 16'h0893;
    16'd24488: out <= 16'hFF4B;    16'd24489: out <= 16'h02BF;    16'd24490: out <= 16'h09B9;    16'd24491: out <= 16'h0515;
    16'd24492: out <= 16'h023B;    16'd24493: out <= 16'h0192;    16'd24494: out <= 16'h0455;    16'd24495: out <= 16'h030B;
    16'd24496: out <= 16'h0225;    16'd24497: out <= 16'h0889;    16'd24498: out <= 16'h065B;    16'd24499: out <= 16'h0A02;
    16'd24500: out <= 16'h011A;    16'd24501: out <= 16'h01D2;    16'd24502: out <= 16'h0879;    16'd24503: out <= 16'h0714;
    16'd24504: out <= 16'h06D1;    16'd24505: out <= 16'h0069;    16'd24506: out <= 16'hFF19;    16'd24507: out <= 16'h028E;
    16'd24508: out <= 16'h0042;    16'd24509: out <= 16'h0826;    16'd24510: out <= 16'hFDF0;    16'd24511: out <= 16'h05B6;
    16'd24512: out <= 16'h0240;    16'd24513: out <= 16'hFAF5;    16'd24514: out <= 16'hFE53;    16'd24515: out <= 16'h0534;
    16'd24516: out <= 16'h0391;    16'd24517: out <= 16'h0403;    16'd24518: out <= 16'h0232;    16'd24519: out <= 16'h08E2;
    16'd24520: out <= 16'h088B;    16'd24521: out <= 16'h0334;    16'd24522: out <= 16'h0946;    16'd24523: out <= 16'hFEF2;
    16'd24524: out <= 16'h0279;    16'd24525: out <= 16'h02EA;    16'd24526: out <= 16'h03EF;    16'd24527: out <= 16'h0EAF;
    16'd24528: out <= 16'h01E6;    16'd24529: out <= 16'h06FB;    16'd24530: out <= 16'h0762;    16'd24531: out <= 16'h07DE;
    16'd24532: out <= 16'h09D8;    16'd24533: out <= 16'h08E4;    16'd24534: out <= 16'h0149;    16'd24535: out <= 16'hFB21;
    16'd24536: out <= 16'h02BB;    16'd24537: out <= 16'h046B;    16'd24538: out <= 16'h034E;    16'd24539: out <= 16'h033C;
    16'd24540: out <= 16'h0A20;    16'd24541: out <= 16'hFD90;    16'd24542: out <= 16'hFE56;    16'd24543: out <= 16'h0694;
    16'd24544: out <= 16'h08B1;    16'd24545: out <= 16'h0079;    16'd24546: out <= 16'hFE69;    16'd24547: out <= 16'hFE87;
    16'd24548: out <= 16'hF707;    16'd24549: out <= 16'h0040;    16'd24550: out <= 16'hF8FB;    16'd24551: out <= 16'hFF30;
    16'd24552: out <= 16'h018D;    16'd24553: out <= 16'h055C;    16'd24554: out <= 16'h002A;    16'd24555: out <= 16'h0122;
    16'd24556: out <= 16'h058B;    16'd24557: out <= 16'hFFE1;    16'd24558: out <= 16'hFEEE;    16'd24559: out <= 16'h05FF;
    16'd24560: out <= 16'h0521;    16'd24561: out <= 16'hFB7C;    16'd24562: out <= 16'h002B;    16'd24563: out <= 16'hFE36;
    16'd24564: out <= 16'h0226;    16'd24565: out <= 16'h004C;    16'd24566: out <= 16'hFC8C;    16'd24567: out <= 16'h0364;
    16'd24568: out <= 16'h02B8;    16'd24569: out <= 16'hF9D9;    16'd24570: out <= 16'h0827;    16'd24571: out <= 16'h0368;
    16'd24572: out <= 16'h04AF;    16'd24573: out <= 16'hFA3A;    16'd24574: out <= 16'hFFA1;    16'd24575: out <= 16'hFE9F;
    16'd24576: out <= 16'h00B7;    16'd24577: out <= 16'h032A;    16'd24578: out <= 16'hFFBF;    16'd24579: out <= 16'h006B;
    16'd24580: out <= 16'hFE66;    16'd24581: out <= 16'hFD66;    16'd24582: out <= 16'h00D2;    16'd24583: out <= 16'h016F;
    16'd24584: out <= 16'h05DE;    16'd24585: out <= 16'h0065;    16'd24586: out <= 16'hFEAE;    16'd24587: out <= 16'hFCAC;
    16'd24588: out <= 16'hFDE5;    16'd24589: out <= 16'h0365;    16'd24590: out <= 16'hFB7D;    16'd24591: out <= 16'h0382;
    16'd24592: out <= 16'h038E;    16'd24593: out <= 16'h0944;    16'd24594: out <= 16'h01EB;    16'd24595: out <= 16'h0390;
    16'd24596: out <= 16'hFB0A;    16'd24597: out <= 16'hF512;    16'd24598: out <= 16'h044C;    16'd24599: out <= 16'h08FC;
    16'd24600: out <= 16'hFC7C;    16'd24601: out <= 16'hFF5D;    16'd24602: out <= 16'hFCBD;    16'd24603: out <= 16'h052B;
    16'd24604: out <= 16'h0021;    16'd24605: out <= 16'h05E4;    16'd24606: out <= 16'h06BE;    16'd24607: out <= 16'h0346;
    16'd24608: out <= 16'h01D4;    16'd24609: out <= 16'h0497;    16'd24610: out <= 16'h0856;    16'd24611: out <= 16'h0398;
    16'd24612: out <= 16'h0379;    16'd24613: out <= 16'h004E;    16'd24614: out <= 16'h09E3;    16'd24615: out <= 16'h0314;
    16'd24616: out <= 16'h05E5;    16'd24617: out <= 16'h05E8;    16'd24618: out <= 16'h0605;    16'd24619: out <= 16'h05E5;
    16'd24620: out <= 16'hFF69;    16'd24621: out <= 16'h08A4;    16'd24622: out <= 16'h02D5;    16'd24623: out <= 16'h0560;
    16'd24624: out <= 16'h038A;    16'd24625: out <= 16'hFCDA;    16'd24626: out <= 16'h074A;    16'd24627: out <= 16'h04C3;
    16'd24628: out <= 16'h0904;    16'd24629: out <= 16'h0240;    16'd24630: out <= 16'h047A;    16'd24631: out <= 16'hFFB7;
    16'd24632: out <= 16'h030B;    16'd24633: out <= 16'h0BB8;    16'd24634: out <= 16'h0683;    16'd24635: out <= 16'h0A67;
    16'd24636: out <= 16'h04FA;    16'd24637: out <= 16'h07B9;    16'd24638: out <= 16'h048C;    16'd24639: out <= 16'h01A5;
    16'd24640: out <= 16'h050F;    16'd24641: out <= 16'h0843;    16'd24642: out <= 16'h03F1;    16'd24643: out <= 16'h0504;
    16'd24644: out <= 16'h015C;    16'd24645: out <= 16'h04B8;    16'd24646: out <= 16'h0A25;    16'd24647: out <= 16'h0060;
    16'd24648: out <= 16'h0511;    16'd24649: out <= 16'h001C;    16'd24650: out <= 16'h06E2;    16'd24651: out <= 16'hFD96;
    16'd24652: out <= 16'h01C1;    16'd24653: out <= 16'h0363;    16'd24654: out <= 16'h047C;    16'd24655: out <= 16'hFF2B;
    16'd24656: out <= 16'hF8C6;    16'd24657: out <= 16'h0560;    16'd24658: out <= 16'hFF15;    16'd24659: out <= 16'h0297;
    16'd24660: out <= 16'h03C1;    16'd24661: out <= 16'h084B;    16'd24662: out <= 16'h071B;    16'd24663: out <= 16'h0A5B;
    16'd24664: out <= 16'h02AE;    16'd24665: out <= 16'h01F1;    16'd24666: out <= 16'hFAF8;    16'd24667: out <= 16'hFB5A;
    16'd24668: out <= 16'h06DC;    16'd24669: out <= 16'h07B1;    16'd24670: out <= 16'hFBDB;    16'd24671: out <= 16'hFB47;
    16'd24672: out <= 16'h05F2;    16'd24673: out <= 16'hFBD7;    16'd24674: out <= 16'hFC66;    16'd24675: out <= 16'h0071;
    16'd24676: out <= 16'hFC6E;    16'd24677: out <= 16'h0212;    16'd24678: out <= 16'h0E26;    16'd24679: out <= 16'h07A5;
    16'd24680: out <= 16'h0481;    16'd24681: out <= 16'h04CD;    16'd24682: out <= 16'hFFBE;    16'd24683: out <= 16'h018F;
    16'd24684: out <= 16'h030F;    16'd24685: out <= 16'h0159;    16'd24686: out <= 16'h0608;    16'd24687: out <= 16'h071F;
    16'd24688: out <= 16'h06BC;    16'd24689: out <= 16'hFC18;    16'd24690: out <= 16'h0382;    16'd24691: out <= 16'h0374;
    16'd24692: out <= 16'h05E0;    16'd24693: out <= 16'h060A;    16'd24694: out <= 16'h03AA;    16'd24695: out <= 16'h00A4;
    16'd24696: out <= 16'h0651;    16'd24697: out <= 16'h0061;    16'd24698: out <= 16'h0217;    16'd24699: out <= 16'h0501;
    16'd24700: out <= 16'hFF38;    16'd24701: out <= 16'hFB7A;    16'd24702: out <= 16'h00AE;    16'd24703: out <= 16'h06EB;
    16'd24704: out <= 16'h02E3;    16'd24705: out <= 16'h0A22;    16'd24706: out <= 16'h06C6;    16'd24707: out <= 16'hFAC2;
    16'd24708: out <= 16'hFE10;    16'd24709: out <= 16'h0061;    16'd24710: out <= 16'h0381;    16'd24711: out <= 16'hFDE7;
    16'd24712: out <= 16'h0325;    16'd24713: out <= 16'h0919;    16'd24714: out <= 16'h050A;    16'd24715: out <= 16'h028C;
    16'd24716: out <= 16'h082C;    16'd24717: out <= 16'h04E3;    16'd24718: out <= 16'h090A;    16'd24719: out <= 16'h00CF;
    16'd24720: out <= 16'h0237;    16'd24721: out <= 16'hFACC;    16'd24722: out <= 16'h0133;    16'd24723: out <= 16'h02DB;
    16'd24724: out <= 16'h0305;    16'd24725: out <= 16'hFDB6;    16'd24726: out <= 16'h0037;    16'd24727: out <= 16'hF938;
    16'd24728: out <= 16'h030C;    16'd24729: out <= 16'h0015;    16'd24730: out <= 16'h0596;    16'd24731: out <= 16'h01D9;
    16'd24732: out <= 16'h053D;    16'd24733: out <= 16'h026C;    16'd24734: out <= 16'h0143;    16'd24735: out <= 16'hFF21;
    16'd24736: out <= 16'hFE51;    16'd24737: out <= 16'h07D7;    16'd24738: out <= 16'h0339;    16'd24739: out <= 16'h020D;
    16'd24740: out <= 16'h02BD;    16'd24741: out <= 16'h06B7;    16'd24742: out <= 16'h078C;    16'd24743: out <= 16'h062B;
    16'd24744: out <= 16'h04A4;    16'd24745: out <= 16'h0108;    16'd24746: out <= 16'hFD67;    16'd24747: out <= 16'h034E;
    16'd24748: out <= 16'h029E;    16'd24749: out <= 16'h02E9;    16'd24750: out <= 16'h0391;    16'd24751: out <= 16'h0075;
    16'd24752: out <= 16'h0861;    16'd24753: out <= 16'hFF2A;    16'd24754: out <= 16'hFF30;    16'd24755: out <= 16'h07EA;
    16'd24756: out <= 16'h010A;    16'd24757: out <= 16'h0B4D;    16'd24758: out <= 16'h00E5;    16'd24759: out <= 16'hFE7E;
    16'd24760: out <= 16'h03BE;    16'd24761: out <= 16'h06F1;    16'd24762: out <= 16'h077D;    16'd24763: out <= 16'h002D;
    16'd24764: out <= 16'h066E;    16'd24765: out <= 16'h00DD;    16'd24766: out <= 16'hFE2C;    16'd24767: out <= 16'h0163;
    16'd24768: out <= 16'h0638;    16'd24769: out <= 16'h069B;    16'd24770: out <= 16'h0545;    16'd24771: out <= 16'h0033;
    16'd24772: out <= 16'h016A;    16'd24773: out <= 16'h025D;    16'd24774: out <= 16'h0741;    16'd24775: out <= 16'hFDA1;
    16'd24776: out <= 16'h079B;    16'd24777: out <= 16'h06FB;    16'd24778: out <= 16'hFB8C;    16'd24779: out <= 16'h0378;
    16'd24780: out <= 16'hF905;    16'd24781: out <= 16'h00DA;    16'd24782: out <= 16'h0246;    16'd24783: out <= 16'hFFAA;
    16'd24784: out <= 16'h06E5;    16'd24785: out <= 16'hFA70;    16'd24786: out <= 16'h00D6;    16'd24787: out <= 16'h04C6;
    16'd24788: out <= 16'h06CB;    16'd24789: out <= 16'h0475;    16'd24790: out <= 16'h0995;    16'd24791: out <= 16'h0C12;
    16'd24792: out <= 16'h0344;    16'd24793: out <= 16'h05B0;    16'd24794: out <= 16'hFF84;    16'd24795: out <= 16'h00DC;
    16'd24796: out <= 16'h03F1;    16'd24797: out <= 16'h05E3;    16'd24798: out <= 16'hFF6E;    16'd24799: out <= 16'h01C7;
    16'd24800: out <= 16'h01B5;    16'd24801: out <= 16'h0247;    16'd24802: out <= 16'h0531;    16'd24803: out <= 16'h020E;
    16'd24804: out <= 16'h0C09;    16'd24805: out <= 16'h0216;    16'd24806: out <= 16'h019B;    16'd24807: out <= 16'hFA4D;
    16'd24808: out <= 16'hFAF1;    16'd24809: out <= 16'hFD8C;    16'd24810: out <= 16'hFB48;    16'd24811: out <= 16'hFECE;
    16'd24812: out <= 16'hFDF6;    16'd24813: out <= 16'h03D4;    16'd24814: out <= 16'hFF9B;    16'd24815: out <= 16'hFD0D;
    16'd24816: out <= 16'hFA72;    16'd24817: out <= 16'hFF01;    16'd24818: out <= 16'hFFD3;    16'd24819: out <= 16'hFFDC;
    16'd24820: out <= 16'hFD08;    16'd24821: out <= 16'hFC72;    16'd24822: out <= 16'h0169;    16'd24823: out <= 16'h00F9;
    16'd24824: out <= 16'h0808;    16'd24825: out <= 16'h00A2;    16'd24826: out <= 16'hFDBE;    16'd24827: out <= 16'h017F;
    16'd24828: out <= 16'hFEFF;    16'd24829: out <= 16'hF882;    16'd24830: out <= 16'hFBC6;    16'd24831: out <= 16'h0595;
    16'd24832: out <= 16'hFB90;    16'd24833: out <= 16'h03A2;    16'd24834: out <= 16'h032A;    16'd24835: out <= 16'hFF09;
    16'd24836: out <= 16'h06BF;    16'd24837: out <= 16'h04F0;    16'd24838: out <= 16'hF97B;    16'd24839: out <= 16'hFFA4;
    16'd24840: out <= 16'hFD1E;    16'd24841: out <= 16'hFFB5;    16'd24842: out <= 16'hF9BC;    16'd24843: out <= 16'h00DB;
    16'd24844: out <= 16'h00D6;    16'd24845: out <= 16'h00C1;    16'd24846: out <= 16'hFFA8;    16'd24847: out <= 16'hFF21;
    16'd24848: out <= 16'h0503;    16'd24849: out <= 16'h07EA;    16'd24850: out <= 16'h0116;    16'd24851: out <= 16'hFF24;
    16'd24852: out <= 16'h000C;    16'd24853: out <= 16'hFF8B;    16'd24854: out <= 16'h03F1;    16'd24855: out <= 16'hFBD3;
    16'd24856: out <= 16'hFC26;    16'd24857: out <= 16'hFEF9;    16'd24858: out <= 16'hFBCD;    16'd24859: out <= 16'h003E;
    16'd24860: out <= 16'h0C16;    16'd24861: out <= 16'h06BC;    16'd24862: out <= 16'h086B;    16'd24863: out <= 16'h05CA;
    16'd24864: out <= 16'h0212;    16'd24865: out <= 16'h0400;    16'd24866: out <= 16'h0D64;    16'd24867: out <= 16'h0659;
    16'd24868: out <= 16'h0397;    16'd24869: out <= 16'hFEFC;    16'd24870: out <= 16'h05A2;    16'd24871: out <= 16'h0D5D;
    16'd24872: out <= 16'h0192;    16'd24873: out <= 16'h01A4;    16'd24874: out <= 16'h01DD;    16'd24875: out <= 16'h07AD;
    16'd24876: out <= 16'h0C8F;    16'd24877: out <= 16'hFE8A;    16'd24878: out <= 16'h08D1;    16'd24879: out <= 16'h01C4;
    16'd24880: out <= 16'h02DF;    16'd24881: out <= 16'h03CA;    16'd24882: out <= 16'hFF14;    16'd24883: out <= 16'h07F5;
    16'd24884: out <= 16'h00C2;    16'd24885: out <= 16'h07F3;    16'd24886: out <= 16'h02EC;    16'd24887: out <= 16'hFE7B;
    16'd24888: out <= 16'hFF03;    16'd24889: out <= 16'h0587;    16'd24890: out <= 16'h02F5;    16'd24891: out <= 16'h06E6;
    16'd24892: out <= 16'h0B3B;    16'd24893: out <= 16'h00F5;    16'd24894: out <= 16'h087D;    16'd24895: out <= 16'h01CF;
    16'd24896: out <= 16'h074B;    16'd24897: out <= 16'h07CB;    16'd24898: out <= 16'hFF8B;    16'd24899: out <= 16'h092C;
    16'd24900: out <= 16'h08D1;    16'd24901: out <= 16'h02D7;    16'd24902: out <= 16'h0898;    16'd24903: out <= 16'h008A;
    16'd24904: out <= 16'h0636;    16'd24905: out <= 16'h06FE;    16'd24906: out <= 16'h01F2;    16'd24907: out <= 16'hFE41;
    16'd24908: out <= 16'h03C6;    16'd24909: out <= 16'h055C;    16'd24910: out <= 16'hF859;    16'd24911: out <= 16'h0247;
    16'd24912: out <= 16'hFDF7;    16'd24913: out <= 16'hFEA3;    16'd24914: out <= 16'h0629;    16'd24915: out <= 16'h0168;
    16'd24916: out <= 16'hFF1D;    16'd24917: out <= 16'hFF3A;    16'd24918: out <= 16'h0501;    16'd24919: out <= 16'h088C;
    16'd24920: out <= 16'h019B;    16'd24921: out <= 16'h0547;    16'd24922: out <= 16'h074A;    16'd24923: out <= 16'h0304;
    16'd24924: out <= 16'h033F;    16'd24925: out <= 16'h0202;    16'd24926: out <= 16'h0609;    16'd24927: out <= 16'hFCC8;
    16'd24928: out <= 16'h011F;    16'd24929: out <= 16'h0045;    16'd24930: out <= 16'h04CC;    16'd24931: out <= 16'hFE97;
    16'd24932: out <= 16'hFC94;    16'd24933: out <= 16'hFDC7;    16'd24934: out <= 16'h046D;    16'd24935: out <= 16'h0C19;
    16'd24936: out <= 16'hF870;    16'd24937: out <= 16'h0675;    16'd24938: out <= 16'h02A3;    16'd24939: out <= 16'h03D2;
    16'd24940: out <= 16'h0118;    16'd24941: out <= 16'h01C9;    16'd24942: out <= 16'hFE1A;    16'd24943: out <= 16'h05C0;
    16'd24944: out <= 16'h08DC;    16'd24945: out <= 16'h02D5;    16'd24946: out <= 16'h06F1;    16'd24947: out <= 16'h045E;
    16'd24948: out <= 16'h036C;    16'd24949: out <= 16'h0BAB;    16'd24950: out <= 16'hFC2A;    16'd24951: out <= 16'h0112;
    16'd24952: out <= 16'h00DF;    16'd24953: out <= 16'h04E2;    16'd24954: out <= 16'h0835;    16'd24955: out <= 16'hFBF7;
    16'd24956: out <= 16'h03C0;    16'd24957: out <= 16'h0701;    16'd24958: out <= 16'h00BD;    16'd24959: out <= 16'h0808;
    16'd24960: out <= 16'h09D8;    16'd24961: out <= 16'hFCB2;    16'd24962: out <= 16'h083C;    16'd24963: out <= 16'h0BEB;
    16'd24964: out <= 16'hFF72;    16'd24965: out <= 16'h019E;    16'd24966: out <= 16'h04DB;    16'd24967: out <= 16'h0877;
    16'd24968: out <= 16'h0025;    16'd24969: out <= 16'hFD1A;    16'd24970: out <= 16'h018C;    16'd24971: out <= 16'h0497;
    16'd24972: out <= 16'h0839;    16'd24973: out <= 16'h041E;    16'd24974: out <= 16'h0276;    16'd24975: out <= 16'h0414;
    16'd24976: out <= 16'h0471;    16'd24977: out <= 16'hFDEE;    16'd24978: out <= 16'hFD4B;    16'd24979: out <= 16'hFC5E;
    16'd24980: out <= 16'h0297;    16'd24981: out <= 16'h05CD;    16'd24982: out <= 16'h03DF;    16'd24983: out <= 16'h059C;
    16'd24984: out <= 16'hFA9D;    16'd24985: out <= 16'h1052;    16'd24986: out <= 16'h06DE;    16'd24987: out <= 16'h0967;
    16'd24988: out <= 16'h05B6;    16'd24989: out <= 16'h099D;    16'd24990: out <= 16'h073F;    16'd24991: out <= 16'h04B6;
    16'd24992: out <= 16'hFFB5;    16'd24993: out <= 16'hFCB7;    16'd24994: out <= 16'h05A5;    16'd24995: out <= 16'h08EA;
    16'd24996: out <= 16'hFF78;    16'd24997: out <= 16'h0A55;    16'd24998: out <= 16'h0A21;    16'd24999: out <= 16'hFF69;
    16'd25000: out <= 16'h013F;    16'd25001: out <= 16'h0032;    16'd25002: out <= 16'h1117;    16'd25003: out <= 16'hFF41;
    16'd25004: out <= 16'h08D5;    16'd25005: out <= 16'h018D;    16'd25006: out <= 16'h0411;    16'd25007: out <= 16'h0600;
    16'd25008: out <= 16'h042B;    16'd25009: out <= 16'h0A73;    16'd25010: out <= 16'hFF75;    16'd25011: out <= 16'h02F5;
    16'd25012: out <= 16'h05A7;    16'd25013: out <= 16'hFF19;    16'd25014: out <= 16'h092E;    16'd25015: out <= 16'h07E9;
    16'd25016: out <= 16'h075D;    16'd25017: out <= 16'h0674;    16'd25018: out <= 16'hFC33;    16'd25019: out <= 16'h0620;
    16'd25020: out <= 16'h065A;    16'd25021: out <= 16'h0699;    16'd25022: out <= 16'h0B32;    16'd25023: out <= 16'h0566;
    16'd25024: out <= 16'h0AF3;    16'd25025: out <= 16'h03AC;    16'd25026: out <= 16'hFD3F;    16'd25027: out <= 16'h01B9;
    16'd25028: out <= 16'hFDBE;    16'd25029: out <= 16'h0523;    16'd25030: out <= 16'h0159;    16'd25031: out <= 16'hFE76;
    16'd25032: out <= 16'h05D7;    16'd25033: out <= 16'h03FA;    16'd25034: out <= 16'h0539;    16'd25035: out <= 16'hFB0F;
    16'd25036: out <= 16'h01FB;    16'd25037: out <= 16'hFFFC;    16'd25038: out <= 16'h045C;    16'd25039: out <= 16'h04C6;
    16'd25040: out <= 16'hFDE7;    16'd25041: out <= 16'h02A2;    16'd25042: out <= 16'h0329;    16'd25043: out <= 16'h02D8;
    16'd25044: out <= 16'h05BA;    16'd25045: out <= 16'h028E;    16'd25046: out <= 16'hFFC9;    16'd25047: out <= 16'h0837;
    16'd25048: out <= 16'hFDBF;    16'd25049: out <= 16'hFE68;    16'd25050: out <= 16'h028C;    16'd25051: out <= 16'h053F;
    16'd25052: out <= 16'h0144;    16'd25053: out <= 16'hFE8C;    16'd25054: out <= 16'h0048;    16'd25055: out <= 16'h0049;
    16'd25056: out <= 16'h011A;    16'd25057: out <= 16'h01CA;    16'd25058: out <= 16'hFBD5;    16'd25059: out <= 16'hFEEE;
    16'd25060: out <= 16'h03CA;    16'd25061: out <= 16'h0568;    16'd25062: out <= 16'hFAC1;    16'd25063: out <= 16'hF835;
    16'd25064: out <= 16'h011F;    16'd25065: out <= 16'hFDC4;    16'd25066: out <= 16'hFB20;    16'd25067: out <= 16'hFB54;
    16'd25068: out <= 16'h02AF;    16'd25069: out <= 16'hFEA1;    16'd25070: out <= 16'hFED7;    16'd25071: out <= 16'hF744;
    16'd25072: out <= 16'h03DB;    16'd25073: out <= 16'h0537;    16'd25074: out <= 16'hFD33;    16'd25075: out <= 16'h040D;
    16'd25076: out <= 16'hFC6A;    16'd25077: out <= 16'h04AC;    16'd25078: out <= 16'hFDEC;    16'd25079: out <= 16'hFAE1;
    16'd25080: out <= 16'hFFA6;    16'd25081: out <= 16'h0690;    16'd25082: out <= 16'h009E;    16'd25083: out <= 16'h0188;
    16'd25084: out <= 16'h035B;    16'd25085: out <= 16'hFC99;    16'd25086: out <= 16'h0472;    16'd25087: out <= 16'hF9EA;
    16'd25088: out <= 16'hFADA;    16'd25089: out <= 16'hFFAC;    16'd25090: out <= 16'hFC53;    16'd25091: out <= 16'h046D;
    16'd25092: out <= 16'hFF52;    16'd25093: out <= 16'h0068;    16'd25094: out <= 16'hFEFB;    16'd25095: out <= 16'hFFC5;
    16'd25096: out <= 16'hF9A5;    16'd25097: out <= 16'hFDA7;    16'd25098: out <= 16'hFFA0;    16'd25099: out <= 16'h045B;
    16'd25100: out <= 16'hFF5F;    16'd25101: out <= 16'h0473;    16'd25102: out <= 16'h03DB;    16'd25103: out <= 16'hF96E;
    16'd25104: out <= 16'h0232;    16'd25105: out <= 16'hFE20;    16'd25106: out <= 16'hF4A7;    16'd25107: out <= 16'hFCC1;
    16'd25108: out <= 16'h0401;    16'd25109: out <= 16'h012F;    16'd25110: out <= 16'hFC77;    16'd25111: out <= 16'hFF72;
    16'd25112: out <= 16'hFE91;    16'd25113: out <= 16'h05E4;    16'd25114: out <= 16'h0171;    16'd25115: out <= 16'h0083;
    16'd25116: out <= 16'h010B;    16'd25117: out <= 16'h01F4;    16'd25118: out <= 16'h05E9;    16'd25119: out <= 16'h019D;
    16'd25120: out <= 16'hFFDC;    16'd25121: out <= 16'h06C5;    16'd25122: out <= 16'h0469;    16'd25123: out <= 16'hFDC8;
    16'd25124: out <= 16'hFE2F;    16'd25125: out <= 16'h03FB;    16'd25126: out <= 16'h0227;    16'd25127: out <= 16'h034E;
    16'd25128: out <= 16'h049D;    16'd25129: out <= 16'hFEBB;    16'd25130: out <= 16'h075F;    16'd25131: out <= 16'h003E;
    16'd25132: out <= 16'h0569;    16'd25133: out <= 16'h0318;    16'd25134: out <= 16'h0471;    16'd25135: out <= 16'h02C7;
    16'd25136: out <= 16'h0725;    16'd25137: out <= 16'h0AE0;    16'd25138: out <= 16'h0395;    16'd25139: out <= 16'h00C2;
    16'd25140: out <= 16'h08F9;    16'd25141: out <= 16'hFF13;    16'd25142: out <= 16'hFE12;    16'd25143: out <= 16'h059F;
    16'd25144: out <= 16'hFF82;    16'd25145: out <= 16'hF94B;    16'd25146: out <= 16'h07F3;    16'd25147: out <= 16'h04A9;
    16'd25148: out <= 16'hFE07;    16'd25149: out <= 16'hFEA5;    16'd25150: out <= 16'h00F8;    16'd25151: out <= 16'hFEC0;
    16'd25152: out <= 16'h0845;    16'd25153: out <= 16'h04F5;    16'd25154: out <= 16'h061A;    16'd25155: out <= 16'h023E;
    16'd25156: out <= 16'h0181;    16'd25157: out <= 16'h0580;    16'd25158: out <= 16'h0246;    16'd25159: out <= 16'hFFD1;
    16'd25160: out <= 16'h017D;    16'd25161: out <= 16'h0102;    16'd25162: out <= 16'h00B4;    16'd25163: out <= 16'h059F;
    16'd25164: out <= 16'h061E;    16'd25165: out <= 16'h0386;    16'd25166: out <= 16'h06E9;    16'd25167: out <= 16'h016F;
    16'd25168: out <= 16'hFE36;    16'd25169: out <= 16'h075C;    16'd25170: out <= 16'h03EF;    16'd25171: out <= 16'h04B0;
    16'd25172: out <= 16'h0339;    16'd25173: out <= 16'hFEFD;    16'd25174: out <= 16'h06EC;    16'd25175: out <= 16'h03AA;
    16'd25176: out <= 16'h08E0;    16'd25177: out <= 16'hFFFF;    16'd25178: out <= 16'h07ED;    16'd25179: out <= 16'hFB0A;
    16'd25180: out <= 16'h040F;    16'd25181: out <= 16'hFE58;    16'd25182: out <= 16'h00F5;    16'd25183: out <= 16'hFF27;
    16'd25184: out <= 16'hFFA8;    16'd25185: out <= 16'h02C9;    16'd25186: out <= 16'h043D;    16'd25187: out <= 16'h05A9;
    16'd25188: out <= 16'h01D1;    16'd25189: out <= 16'h0143;    16'd25190: out <= 16'h00B1;    16'd25191: out <= 16'h062A;
    16'd25192: out <= 16'hFF72;    16'd25193: out <= 16'h05B7;    16'd25194: out <= 16'h00AD;    16'd25195: out <= 16'h05AB;
    16'd25196: out <= 16'h0353;    16'd25197: out <= 16'h03A5;    16'd25198: out <= 16'h0613;    16'd25199: out <= 16'h03C0;
    16'd25200: out <= 16'h0316;    16'd25201: out <= 16'h0BD1;    16'd25202: out <= 16'h093F;    16'd25203: out <= 16'h03A9;
    16'd25204: out <= 16'h0274;    16'd25205: out <= 16'h0589;    16'd25206: out <= 16'h00C0;    16'd25207: out <= 16'hFFFB;
    16'd25208: out <= 16'h0651;    16'd25209: out <= 16'h0597;    16'd25210: out <= 16'h009E;    16'd25211: out <= 16'h08E7;
    16'd25212: out <= 16'h009C;    16'd25213: out <= 16'h0521;    16'd25214: out <= 16'hFF73;    16'd25215: out <= 16'h01F0;
    16'd25216: out <= 16'h0AB0;    16'd25217: out <= 16'h0B7B;    16'd25218: out <= 16'hFBBC;    16'd25219: out <= 16'h0B42;
    16'd25220: out <= 16'h02EB;    16'd25221: out <= 16'h001B;    16'd25222: out <= 16'h0481;    16'd25223: out <= 16'h08D3;
    16'd25224: out <= 16'hFC47;    16'd25225: out <= 16'h00D1;    16'd25226: out <= 16'h0533;    16'd25227: out <= 16'hFC4A;
    16'd25228: out <= 16'h0411;    16'd25229: out <= 16'h04C1;    16'd25230: out <= 16'hFB37;    16'd25231: out <= 16'hFE49;
    16'd25232: out <= 16'hFCB4;    16'd25233: out <= 16'hFF33;    16'd25234: out <= 16'h0250;    16'd25235: out <= 16'hFD00;
    16'd25236: out <= 16'hFEE0;    16'd25237: out <= 16'h07CC;    16'd25238: out <= 16'h0637;    16'd25239: out <= 16'h0B20;
    16'd25240: out <= 16'hFBF0;    16'd25241: out <= 16'h0680;    16'd25242: out <= 16'h0254;    16'd25243: out <= 16'h0190;
    16'd25244: out <= 16'h0441;    16'd25245: out <= 16'h04F0;    16'd25246: out <= 16'hFBCA;    16'd25247: out <= 16'h0471;
    16'd25248: out <= 16'h0200;    16'd25249: out <= 16'h0990;    16'd25250: out <= 16'h0749;    16'd25251: out <= 16'hFF95;
    16'd25252: out <= 16'hFF8E;    16'd25253: out <= 16'h04BD;    16'd25254: out <= 16'h042F;    16'd25255: out <= 16'h0253;
    16'd25256: out <= 16'h0287;    16'd25257: out <= 16'h0063;    16'd25258: out <= 16'h00C5;    16'd25259: out <= 16'h00EC;
    16'd25260: out <= 16'hFDFB;    16'd25261: out <= 16'h042B;    16'd25262: out <= 16'h0930;    16'd25263: out <= 16'h0215;
    16'd25264: out <= 16'hFA77;    16'd25265: out <= 16'h039B;    16'd25266: out <= 16'hFEBB;    16'd25267: out <= 16'h00DE;
    16'd25268: out <= 16'h0362;    16'd25269: out <= 16'hFDFC;    16'd25270: out <= 16'h06EA;    16'd25271: out <= 16'h00DD;
    16'd25272: out <= 16'h0005;    16'd25273: out <= 16'h0239;    16'd25274: out <= 16'h016F;    16'd25275: out <= 16'h034C;
    16'd25276: out <= 16'h0390;    16'd25277: out <= 16'h0513;    16'd25278: out <= 16'h07FA;    16'd25279: out <= 16'h01B0;
    16'd25280: out <= 16'h03E3;    16'd25281: out <= 16'h020E;    16'd25282: out <= 16'h054E;    16'd25283: out <= 16'h06BF;
    16'd25284: out <= 16'h0163;    16'd25285: out <= 16'h0A70;    16'd25286: out <= 16'hFEDF;    16'd25287: out <= 16'h05CE;
    16'd25288: out <= 16'h0441;    16'd25289: out <= 16'h08A7;    16'd25290: out <= 16'h086F;    16'd25291: out <= 16'h026C;
    16'd25292: out <= 16'h015C;    16'd25293: out <= 16'h01F0;    16'd25294: out <= 16'h052D;    16'd25295: out <= 16'h07C5;
    16'd25296: out <= 16'h00EF;    16'd25297: out <= 16'h0096;    16'd25298: out <= 16'h091D;    16'd25299: out <= 16'h080E;
    16'd25300: out <= 16'h0276;    16'd25301: out <= 16'h0759;    16'd25302: out <= 16'h02C1;    16'd25303: out <= 16'h055F;
    16'd25304: out <= 16'h00F3;    16'd25305: out <= 16'h0794;    16'd25306: out <= 16'h015E;    16'd25307: out <= 16'h0B0E;
    16'd25308: out <= 16'h0173;    16'd25309: out <= 16'h0658;    16'd25310: out <= 16'hFB3A;    16'd25311: out <= 16'h0313;
    16'd25312: out <= 16'h0296;    16'd25313: out <= 16'h0042;    16'd25314: out <= 16'h02AE;    16'd25315: out <= 16'h017A;
    16'd25316: out <= 16'hFEF7;    16'd25317: out <= 16'h01EA;    16'd25318: out <= 16'h00DE;    16'd25319: out <= 16'hFFD0;
    16'd25320: out <= 16'h0032;    16'd25321: out <= 16'hFE67;    16'd25322: out <= 16'h07E2;    16'd25323: out <= 16'h05E3;
    16'd25324: out <= 16'hFEA5;    16'd25325: out <= 16'hF99F;    16'd25326: out <= 16'h012F;    16'd25327: out <= 16'h0107;
    16'd25328: out <= 16'h03E0;    16'd25329: out <= 16'hFE20;    16'd25330: out <= 16'h006F;    16'd25331: out <= 16'h01A6;
    16'd25332: out <= 16'hFDD8;    16'd25333: out <= 16'hFD96;    16'd25334: out <= 16'h0456;    16'd25335: out <= 16'hFBEC;
    16'd25336: out <= 16'hFE56;    16'd25337: out <= 16'h054A;    16'd25338: out <= 16'hFBFE;    16'd25339: out <= 16'h0385;
    16'd25340: out <= 16'hFB3E;    16'd25341: out <= 16'hFE1F;    16'd25342: out <= 16'hFF0A;    16'd25343: out <= 16'h031E;
    16'd25344: out <= 16'hFF69;    16'd25345: out <= 16'h0245;    16'd25346: out <= 16'h0159;    16'd25347: out <= 16'h0164;
    16'd25348: out <= 16'h05AE;    16'd25349: out <= 16'hFB9E;    16'd25350: out <= 16'hFE67;    16'd25351: out <= 16'hFC6F;
    16'd25352: out <= 16'h0225;    16'd25353: out <= 16'hFE2D;    16'd25354: out <= 16'hFFA8;    16'd25355: out <= 16'h0326;
    16'd25356: out <= 16'hFDE8;    16'd25357: out <= 16'hFF4E;    16'd25358: out <= 16'hFF27;    16'd25359: out <= 16'h0027;
    16'd25360: out <= 16'hFFBA;    16'd25361: out <= 16'h005E;    16'd25362: out <= 16'h00D0;    16'd25363: out <= 16'hFA41;
    16'd25364: out <= 16'hFC63;    16'd25365: out <= 16'hFD0E;    16'd25366: out <= 16'hFF70;    16'd25367: out <= 16'hFB81;
    16'd25368: out <= 16'h015B;    16'd25369: out <= 16'hF9EB;    16'd25370: out <= 16'h01BB;    16'd25371: out <= 16'hFE44;
    16'd25372: out <= 16'h016E;    16'd25373: out <= 16'h0C8A;    16'd25374: out <= 16'h01B4;    16'd25375: out <= 16'h01EC;
    16'd25376: out <= 16'h01DD;    16'd25377: out <= 16'h0178;    16'd25378: out <= 16'h022B;    16'd25379: out <= 16'h0615;
    16'd25380: out <= 16'h06D3;    16'd25381: out <= 16'hFFBA;    16'd25382: out <= 16'h0EAF;    16'd25383: out <= 16'h0AC6;
    16'd25384: out <= 16'h0747;    16'd25385: out <= 16'h0446;    16'd25386: out <= 16'h041A;    16'd25387: out <= 16'h09D9;
    16'd25388: out <= 16'h022B;    16'd25389: out <= 16'h0848;    16'd25390: out <= 16'h0497;    16'd25391: out <= 16'h06C6;
    16'd25392: out <= 16'h0880;    16'd25393: out <= 16'h05DF;    16'd25394: out <= 16'h0774;    16'd25395: out <= 16'h0697;
    16'd25396: out <= 16'h0983;    16'd25397: out <= 16'h0694;    16'd25398: out <= 16'h0168;    16'd25399: out <= 16'h046A;
    16'd25400: out <= 16'hFD92;    16'd25401: out <= 16'h03CD;    16'd25402: out <= 16'h0A4D;    16'd25403: out <= 16'h0909;
    16'd25404: out <= 16'h02DE;    16'd25405: out <= 16'h0481;    16'd25406: out <= 16'h03AE;    16'd25407: out <= 16'h0290;
    16'd25408: out <= 16'h0674;    16'd25409: out <= 16'h05BF;    16'd25410: out <= 16'h05B5;    16'd25411: out <= 16'h0467;
    16'd25412: out <= 16'h008F;    16'd25413: out <= 16'h079F;    16'd25414: out <= 16'hFE8D;    16'd25415: out <= 16'h0263;
    16'd25416: out <= 16'h0054;    16'd25417: out <= 16'hFF36;    16'd25418: out <= 16'hFD32;    16'd25419: out <= 16'h00E1;
    16'd25420: out <= 16'h017D;    16'd25421: out <= 16'h04CA;    16'd25422: out <= 16'h01A6;    16'd25423: out <= 16'h00EE;
    16'd25424: out <= 16'hFAD3;    16'd25425: out <= 16'hFE78;    16'd25426: out <= 16'hFCB8;    16'd25427: out <= 16'hF857;
    16'd25428: out <= 16'h087A;    16'd25429: out <= 16'h02A5;    16'd25430: out <= 16'h0534;    16'd25431: out <= 16'h07E7;
    16'd25432: out <= 16'hFDDD;    16'd25433: out <= 16'h058A;    16'd25434: out <= 16'h031F;    16'd25435: out <= 16'hFB8A;
    16'd25436: out <= 16'hFDD5;    16'd25437: out <= 16'h0103;    16'd25438: out <= 16'h04CC;    16'd25439: out <= 16'h005C;
    16'd25440: out <= 16'h0709;    16'd25441: out <= 16'h0075;    16'd25442: out <= 16'h04B0;    16'd25443: out <= 16'h012B;
    16'd25444: out <= 16'h08A7;    16'd25445: out <= 16'hFD5A;    16'd25446: out <= 16'hF9D3;    16'd25447: out <= 16'h042B;
    16'd25448: out <= 16'h02B6;    16'd25449: out <= 16'h079B;    16'd25450: out <= 16'h0184;    16'd25451: out <= 16'h0318;
    16'd25452: out <= 16'h0654;    16'd25453: out <= 16'hFFF6;    16'd25454: out <= 16'h06D0;    16'd25455: out <= 16'h0743;
    16'd25456: out <= 16'h035A;    16'd25457: out <= 16'h0471;    16'd25458: out <= 16'h0351;    16'd25459: out <= 16'h0423;
    16'd25460: out <= 16'h069F;    16'd25461: out <= 16'h08AD;    16'd25462: out <= 16'h000A;    16'd25463: out <= 16'h055D;
    16'd25464: out <= 16'hFF38;    16'd25465: out <= 16'hFE30;    16'd25466: out <= 16'h01E1;    16'd25467: out <= 16'h03CF;
    16'd25468: out <= 16'h0648;    16'd25469: out <= 16'h0655;    16'd25470: out <= 16'h0386;    16'd25471: out <= 16'h078B;
    16'd25472: out <= 16'h0197;    16'd25473: out <= 16'h040B;    16'd25474: out <= 16'hFF3D;    16'd25475: out <= 16'h0276;
    16'd25476: out <= 16'h00C8;    16'd25477: out <= 16'h0610;    16'd25478: out <= 16'h015A;    16'd25479: out <= 16'h035D;
    16'd25480: out <= 16'h068F;    16'd25481: out <= 16'h07F7;    16'd25482: out <= 16'h0797;    16'd25483: out <= 16'h04EC;
    16'd25484: out <= 16'h06E6;    16'd25485: out <= 16'h035A;    16'd25486: out <= 16'hFA69;    16'd25487: out <= 16'h0D2E;
    16'd25488: out <= 16'h0460;    16'd25489: out <= 16'hFD92;    16'd25490: out <= 16'h036E;    16'd25491: out <= 16'h0041;
    16'd25492: out <= 16'h0AF4;    16'd25493: out <= 16'h0627;    16'd25494: out <= 16'h088A;    16'd25495: out <= 16'hFE95;
    16'd25496: out <= 16'hFF3A;    16'd25497: out <= 16'h0188;    16'd25498: out <= 16'h0422;    16'd25499: out <= 16'h0424;
    16'd25500: out <= 16'h0652;    16'd25501: out <= 16'h0640;    16'd25502: out <= 16'h07FF;    16'd25503: out <= 16'hFEC1;
    16'd25504: out <= 16'h080E;    16'd25505: out <= 16'hFE89;    16'd25506: out <= 16'h02F8;    16'd25507: out <= 16'hFCA9;
    16'd25508: out <= 16'hFFB2;    16'd25509: out <= 16'h009C;    16'd25510: out <= 16'hF911;    16'd25511: out <= 16'hFFCF;
    16'd25512: out <= 16'hFF71;    16'd25513: out <= 16'h011A;    16'd25514: out <= 16'hFDF2;    16'd25515: out <= 16'h067A;
    16'd25516: out <= 16'h0770;    16'd25517: out <= 16'h074A;    16'd25518: out <= 16'h085C;    16'd25519: out <= 16'h05E1;
    16'd25520: out <= 16'h0769;    16'd25521: out <= 16'h05B7;    16'd25522: out <= 16'h00F9;    16'd25523: out <= 16'hF734;
    16'd25524: out <= 16'h0D89;    16'd25525: out <= 16'h04B2;    16'd25526: out <= 16'h01F0;    16'd25527: out <= 16'h043F;
    16'd25528: out <= 16'h04D1;    16'd25529: out <= 16'h04DA;    16'd25530: out <= 16'h0114;    16'd25531: out <= 16'h0564;
    16'd25532: out <= 16'h0681;    16'd25533: out <= 16'h06FA;    16'd25534: out <= 16'h00E3;    16'd25535: out <= 16'h00F3;
    16'd25536: out <= 16'h04BC;    16'd25537: out <= 16'h0779;    16'd25538: out <= 16'h03E8;    16'd25539: out <= 16'h0324;
    16'd25540: out <= 16'hFBEB;    16'd25541: out <= 16'hFA44;    16'd25542: out <= 16'hFEA8;    16'd25543: out <= 16'h08AB;
    16'd25544: out <= 16'h06E7;    16'd25545: out <= 16'h0984;    16'd25546: out <= 16'hFC21;    16'd25547: out <= 16'h0321;
    16'd25548: out <= 16'hFEA7;    16'd25549: out <= 16'h01FD;    16'd25550: out <= 16'h08BE;    16'd25551: out <= 16'h0B62;
    16'd25552: out <= 16'h0386;    16'd25553: out <= 16'h0939;    16'd25554: out <= 16'h01C6;    16'd25555: out <= 16'hFCFB;
    16'd25556: out <= 16'h0024;    16'd25557: out <= 16'h04F2;    16'd25558: out <= 16'hFFC5;    16'd25559: out <= 16'h024D;
    16'd25560: out <= 16'h04ED;    16'd25561: out <= 16'h0796;    16'd25562: out <= 16'h02FA;    16'd25563: out <= 16'h018D;
    16'd25564: out <= 16'h02A5;    16'd25565: out <= 16'hFF33;    16'd25566: out <= 16'h07C6;    16'd25567: out <= 16'hFDF4;
    16'd25568: out <= 16'h0281;    16'd25569: out <= 16'hF9BB;    16'd25570: out <= 16'h03F5;    16'd25571: out <= 16'h06A0;
    16'd25572: out <= 16'h046E;    16'd25573: out <= 16'h04C0;    16'd25574: out <= 16'h03AE;    16'd25575: out <= 16'hFAD9;
    16'd25576: out <= 16'h0236;    16'd25577: out <= 16'hFBAC;    16'd25578: out <= 16'hFD56;    16'd25579: out <= 16'h063C;
    16'd25580: out <= 16'h03E7;    16'd25581: out <= 16'hFA05;    16'd25582: out <= 16'hFF7B;    16'd25583: out <= 16'hFD5A;
    16'd25584: out <= 16'hFF09;    16'd25585: out <= 16'hF964;    16'd25586: out <= 16'h0600;    16'd25587: out <= 16'hFBF5;
    16'd25588: out <= 16'hF96A;    16'd25589: out <= 16'h0289;    16'd25590: out <= 16'h006C;    16'd25591: out <= 16'hFD5C;
    16'd25592: out <= 16'h01E5;    16'd25593: out <= 16'hFF82;    16'd25594: out <= 16'h000C;    16'd25595: out <= 16'h04AB;
    16'd25596: out <= 16'h0556;    16'd25597: out <= 16'hFD32;    16'd25598: out <= 16'hFEED;    16'd25599: out <= 16'h039B;
    16'd25600: out <= 16'h0270;    16'd25601: out <= 16'hFF66;    16'd25602: out <= 16'h02CC;    16'd25603: out <= 16'hFC12;
    16'd25604: out <= 16'hFB80;    16'd25605: out <= 16'h0404;    16'd25606: out <= 16'h0722;    16'd25607: out <= 16'h0184;
    16'd25608: out <= 16'h02D2;    16'd25609: out <= 16'h01FE;    16'd25610: out <= 16'h04C9;    16'd25611: out <= 16'h0295;
    16'd25612: out <= 16'h0779;    16'd25613: out <= 16'hFF52;    16'd25614: out <= 16'hF777;    16'd25615: out <= 16'h00C4;
    16'd25616: out <= 16'hFE03;    16'd25617: out <= 16'h0087;    16'd25618: out <= 16'h07ED;    16'd25619: out <= 16'hFFF9;
    16'd25620: out <= 16'hFE6D;    16'd25621: out <= 16'h0146;    16'd25622: out <= 16'h0184;    16'd25623: out <= 16'hFA9A;
    16'd25624: out <= 16'h02AC;    16'd25625: out <= 16'h0515;    16'd25626: out <= 16'h0533;    16'd25627: out <= 16'h00D7;
    16'd25628: out <= 16'h0428;    16'd25629: out <= 16'h0932;    16'd25630: out <= 16'hFD2E;    16'd25631: out <= 16'hFD51;
    16'd25632: out <= 16'h087B;    16'd25633: out <= 16'hFE22;    16'd25634: out <= 16'h0129;    16'd25635: out <= 16'h09FB;
    16'd25636: out <= 16'h0201;    16'd25637: out <= 16'hFED6;    16'd25638: out <= 16'h01C3;    16'd25639: out <= 16'h059A;
    16'd25640: out <= 16'h0595;    16'd25641: out <= 16'h0245;    16'd25642: out <= 16'h013B;    16'd25643: out <= 16'hFD0D;
    16'd25644: out <= 16'h036E;    16'd25645: out <= 16'h00BC;    16'd25646: out <= 16'h011D;    16'd25647: out <= 16'h0710;
    16'd25648: out <= 16'h0356;    16'd25649: out <= 16'h0BBB;    16'd25650: out <= 16'h0274;    16'd25651: out <= 16'h0217;
    16'd25652: out <= 16'h01A3;    16'd25653: out <= 16'h02D3;    16'd25654: out <= 16'h05D5;    16'd25655: out <= 16'h0109;
    16'd25656: out <= 16'h01EF;    16'd25657: out <= 16'h0704;    16'd25658: out <= 16'h0242;    16'd25659: out <= 16'h0444;
    16'd25660: out <= 16'h08F7;    16'd25661: out <= 16'h08D8;    16'd25662: out <= 16'h0C70;    16'd25663: out <= 16'h00B7;
    16'd25664: out <= 16'h0279;    16'd25665: out <= 16'h02EA;    16'd25666: out <= 16'h0049;    16'd25667: out <= 16'h0211;
    16'd25668: out <= 16'hFDEA;    16'd25669: out <= 16'h0900;    16'd25670: out <= 16'h0843;    16'd25671: out <= 16'h0255;
    16'd25672: out <= 16'h0095;    16'd25673: out <= 16'h0930;    16'd25674: out <= 16'hFB3D;    16'd25675: out <= 16'h02F3;
    16'd25676: out <= 16'h00F1;    16'd25677: out <= 16'hFA41;    16'd25678: out <= 16'h0394;    16'd25679: out <= 16'h0468;
    16'd25680: out <= 16'h016A;    16'd25681: out <= 16'h05F7;    16'd25682: out <= 16'h096C;    16'd25683: out <= 16'h02DC;
    16'd25684: out <= 16'h04EE;    16'd25685: out <= 16'h008F;    16'd25686: out <= 16'h076C;    16'd25687: out <= 16'h02A1;
    16'd25688: out <= 16'hFE07;    16'd25689: out <= 16'h012C;    16'd25690: out <= 16'h0022;    16'd25691: out <= 16'h0117;
    16'd25692: out <= 16'h05F0;    16'd25693: out <= 16'h00FF;    16'd25694: out <= 16'hF8FA;    16'd25695: out <= 16'hF941;
    16'd25696: out <= 16'hFFA0;    16'd25697: out <= 16'hFBCA;    16'd25698: out <= 16'h04F5;    16'd25699: out <= 16'hFFAF;
    16'd25700: out <= 16'hFEB1;    16'd25701: out <= 16'h05B7;    16'd25702: out <= 16'hFDEC;    16'd25703: out <= 16'h0575;
    16'd25704: out <= 16'h0394;    16'd25705: out <= 16'h0B52;    16'd25706: out <= 16'h016A;    16'd25707: out <= 16'hFE1D;
    16'd25708: out <= 16'h0893;    16'd25709: out <= 16'h0A27;    16'd25710: out <= 16'h04D6;    16'd25711: out <= 16'hFE6D;
    16'd25712: out <= 16'hFD82;    16'd25713: out <= 16'h0E8B;    16'd25714: out <= 16'h0795;    16'd25715: out <= 16'hFB94;
    16'd25716: out <= 16'h0128;    16'd25717: out <= 16'h0229;    16'd25718: out <= 16'h0868;    16'd25719: out <= 16'h035A;
    16'd25720: out <= 16'h0718;    16'd25721: out <= 16'h072D;    16'd25722: out <= 16'h01FE;    16'd25723: out <= 16'h07D7;
    16'd25724: out <= 16'h02BB;    16'd25725: out <= 16'h0252;    16'd25726: out <= 16'h005D;    16'd25727: out <= 16'h0734;
    16'd25728: out <= 16'hFFDA;    16'd25729: out <= 16'h028A;    16'd25730: out <= 16'h02A5;    16'd25731: out <= 16'h01F2;
    16'd25732: out <= 16'h009C;    16'd25733: out <= 16'h07DE;    16'd25734: out <= 16'h014C;    16'd25735: out <= 16'h091A;
    16'd25736: out <= 16'h03CC;    16'd25737: out <= 16'h04DE;    16'd25738: out <= 16'h011F;    16'd25739: out <= 16'h03BA;
    16'd25740: out <= 16'h016A;    16'd25741: out <= 16'h0097;    16'd25742: out <= 16'h03CF;    16'd25743: out <= 16'h07FB;
    16'd25744: out <= 16'h024E;    16'd25745: out <= 16'h0697;    16'd25746: out <= 16'h0D4B;    16'd25747: out <= 16'h05C9;
    16'd25748: out <= 16'hFF73;    16'd25749: out <= 16'h067C;    16'd25750: out <= 16'h0423;    16'd25751: out <= 16'hFA3E;
    16'd25752: out <= 16'h0377;    16'd25753: out <= 16'h0387;    16'd25754: out <= 16'h0413;    16'd25755: out <= 16'h060B;
    16'd25756: out <= 16'h0576;    16'd25757: out <= 16'h051C;    16'd25758: out <= 16'h02C1;    16'd25759: out <= 16'h033A;
    16'd25760: out <= 16'h046C;    16'd25761: out <= 16'h0324;    16'd25762: out <= 16'h0005;    16'd25763: out <= 16'hFB77;
    16'd25764: out <= 16'h009E;    16'd25765: out <= 16'hFF98;    16'd25766: out <= 16'h084C;    16'd25767: out <= 16'h0176;
    16'd25768: out <= 16'hFCBA;    16'd25769: out <= 16'h0345;    16'd25770: out <= 16'hFD84;    16'd25771: out <= 16'h02B3;
    16'd25772: out <= 16'h01F0;    16'd25773: out <= 16'hF9B6;    16'd25774: out <= 16'h07FE;    16'd25775: out <= 16'h0510;
    16'd25776: out <= 16'h02C8;    16'd25777: out <= 16'h0165;    16'd25778: out <= 16'h028A;    16'd25779: out <= 16'h0307;
    16'd25780: out <= 16'hFCE3;    16'd25781: out <= 16'hFE2E;    16'd25782: out <= 16'h09C5;    16'd25783: out <= 16'h034B;
    16'd25784: out <= 16'h0293;    16'd25785: out <= 16'h02BF;    16'd25786: out <= 16'hFB6B;    16'd25787: out <= 16'h04FC;
    16'd25788: out <= 16'hFC95;    16'd25789: out <= 16'hFD7D;    16'd25790: out <= 16'h09D9;    16'd25791: out <= 16'h032B;
    16'd25792: out <= 16'h043A;    16'd25793: out <= 16'hFC8C;    16'd25794: out <= 16'h083C;    16'd25795: out <= 16'h0281;
    16'd25796: out <= 16'h01A5;    16'd25797: out <= 16'h0406;    16'd25798: out <= 16'hFFC0;    16'd25799: out <= 16'h0274;
    16'd25800: out <= 16'h03DC;    16'd25801: out <= 16'h0083;    16'd25802: out <= 16'h05A6;    16'd25803: out <= 16'h059A;
    16'd25804: out <= 16'h014E;    16'd25805: out <= 16'h097A;    16'd25806: out <= 16'hFF40;    16'd25807: out <= 16'h05E6;
    16'd25808: out <= 16'hFECE;    16'd25809: out <= 16'h040C;    16'd25810: out <= 16'h098B;    16'd25811: out <= 16'h05A6;
    16'd25812: out <= 16'h01E5;    16'd25813: out <= 16'h0566;    16'd25814: out <= 16'h0755;    16'd25815: out <= 16'h00EB;
    16'd25816: out <= 16'h011E;    16'd25817: out <= 16'h066E;    16'd25818: out <= 16'h06A2;    16'd25819: out <= 16'h0960;
    16'd25820: out <= 16'hFFB7;    16'd25821: out <= 16'hF825;    16'd25822: out <= 16'h0296;    16'd25823: out <= 16'h0272;
    16'd25824: out <= 16'hF7B9;    16'd25825: out <= 16'hFC1E;    16'd25826: out <= 16'hFF68;    16'd25827: out <= 16'h0304;
    16'd25828: out <= 16'h038E;    16'd25829: out <= 16'h0271;    16'd25830: out <= 16'h0222;    16'd25831: out <= 16'hFB45;
    16'd25832: out <= 16'h04DD;    16'd25833: out <= 16'hFB93;    16'd25834: out <= 16'hFA80;    16'd25835: out <= 16'hFA95;
    16'd25836: out <= 16'h00E2;    16'd25837: out <= 16'hFF07;    16'd25838: out <= 16'hFAD0;    16'd25839: out <= 16'hFE99;
    16'd25840: out <= 16'hFDB6;    16'd25841: out <= 16'h030F;    16'd25842: out <= 16'hFCFE;    16'd25843: out <= 16'h07AC;
    16'd25844: out <= 16'hFC5B;    16'd25845: out <= 16'h00A7;    16'd25846: out <= 16'h0448;    16'd25847: out <= 16'hFA41;
    16'd25848: out <= 16'hFC22;    16'd25849: out <= 16'h02E1;    16'd25850: out <= 16'hFE66;    16'd25851: out <= 16'h08FD;
    16'd25852: out <= 16'h0320;    16'd25853: out <= 16'h0548;    16'd25854: out <= 16'hFC94;    16'd25855: out <= 16'h03A5;
    16'd25856: out <= 16'hFDCD;    16'd25857: out <= 16'hFEE5;    16'd25858: out <= 16'h0013;    16'd25859: out <= 16'hFEE1;
    16'd25860: out <= 16'h0148;    16'd25861: out <= 16'h0135;    16'd25862: out <= 16'hFB16;    16'd25863: out <= 16'hFB17;
    16'd25864: out <= 16'h0244;    16'd25865: out <= 16'hFEF2;    16'd25866: out <= 16'h013D;    16'd25867: out <= 16'hFD6E;
    16'd25868: out <= 16'hFB76;    16'd25869: out <= 16'hF9F9;    16'd25870: out <= 16'h0394;    16'd25871: out <= 16'h007C;
    16'd25872: out <= 16'h0164;    16'd25873: out <= 16'h0403;    16'd25874: out <= 16'h0134;    16'd25875: out <= 16'h041B;
    16'd25876: out <= 16'hFD8F;    16'd25877: out <= 16'hFBDD;    16'd25878: out <= 16'h096B;    16'd25879: out <= 16'hFFEB;
    16'd25880: out <= 16'h0179;    16'd25881: out <= 16'h0078;    16'd25882: out <= 16'hFAE8;    16'd25883: out <= 16'hFBDD;
    16'd25884: out <= 16'hF8A0;    16'd25885: out <= 16'hFE8E;    16'd25886: out <= 16'h0501;    16'd25887: out <= 16'hFEA7;
    16'd25888: out <= 16'h0185;    16'd25889: out <= 16'h0730;    16'd25890: out <= 16'h04EB;    16'd25891: out <= 16'h0615;
    16'd25892: out <= 16'h0187;    16'd25893: out <= 16'h0268;    16'd25894: out <= 16'h0827;    16'd25895: out <= 16'h088C;
    16'd25896: out <= 16'h0468;    16'd25897: out <= 16'h0446;    16'd25898: out <= 16'hFF27;    16'd25899: out <= 16'h0485;
    16'd25900: out <= 16'hFCD5;    16'd25901: out <= 16'h0329;    16'd25902: out <= 16'hFE0B;    16'd25903: out <= 16'hFEFF;
    16'd25904: out <= 16'h0180;    16'd25905: out <= 16'hFEBC;    16'd25906: out <= 16'hFEBB;    16'd25907: out <= 16'h0682;
    16'd25908: out <= 16'h0217;    16'd25909: out <= 16'h0102;    16'd25910: out <= 16'h07EE;    16'd25911: out <= 16'hFEEE;
    16'd25912: out <= 16'h0589;    16'd25913: out <= 16'h006A;    16'd25914: out <= 16'h02E0;    16'd25915: out <= 16'hFFE3;
    16'd25916: out <= 16'h0997;    16'd25917: out <= 16'hFFD3;    16'd25918: out <= 16'h0198;    16'd25919: out <= 16'h0A84;
    16'd25920: out <= 16'h005F;    16'd25921: out <= 16'h0EE6;    16'd25922: out <= 16'hFA2C;    16'd25923: out <= 16'h0274;
    16'd25924: out <= 16'h00E3;    16'd25925: out <= 16'h006D;    16'd25926: out <= 16'h0452;    16'd25927: out <= 16'hFF0D;
    16'd25928: out <= 16'h04FF;    16'd25929: out <= 16'h07C9;    16'd25930: out <= 16'hFEEF;    16'd25931: out <= 16'h02AB;
    16'd25932: out <= 16'h04D0;    16'd25933: out <= 16'hFE52;    16'd25934: out <= 16'h04B3;    16'd25935: out <= 16'h010C;
    16'd25936: out <= 16'h051D;    16'd25937: out <= 16'h0564;    16'd25938: out <= 16'hFE67;    16'd25939: out <= 16'h0348;
    16'd25940: out <= 16'h06BA;    16'd25941: out <= 16'h03E1;    16'd25942: out <= 16'h06E1;    16'd25943: out <= 16'h0946;
    16'd25944: out <= 16'hFE0B;    16'd25945: out <= 16'h04C2;    16'd25946: out <= 16'h0701;    16'd25947: out <= 16'h08E6;
    16'd25948: out <= 16'hFBFE;    16'd25949: out <= 16'hFF48;    16'd25950: out <= 16'h02BF;    16'd25951: out <= 16'hF6D9;
    16'd25952: out <= 16'hFD1C;    16'd25953: out <= 16'hF97D;    16'd25954: out <= 16'hF9F3;    16'd25955: out <= 16'h0306;
    16'd25956: out <= 16'h00B9;    16'd25957: out <= 16'hFE8B;    16'd25958: out <= 16'h082A;    16'd25959: out <= 16'h0C20;
    16'd25960: out <= 16'h0492;    16'd25961: out <= 16'h0100;    16'd25962: out <= 16'h042F;    16'd25963: out <= 16'h0151;
    16'd25964: out <= 16'h01D9;    16'd25965: out <= 16'hFF27;    16'd25966: out <= 16'h0A21;    16'd25967: out <= 16'hFEA7;
    16'd25968: out <= 16'h0181;    16'd25969: out <= 16'h0997;    16'd25970: out <= 16'h06FB;    16'd25971: out <= 16'h00B3;
    16'd25972: out <= 16'h045F;    16'd25973: out <= 16'h0817;    16'd25974: out <= 16'h060B;    16'd25975: out <= 16'hFF9E;
    16'd25976: out <= 16'h0537;    16'd25977: out <= 16'hFFB7;    16'd25978: out <= 16'h0586;    16'd25979: out <= 16'hFE74;
    16'd25980: out <= 16'h0321;    16'd25981: out <= 16'h0685;    16'd25982: out <= 16'hFE2C;    16'd25983: out <= 16'h07F5;
    16'd25984: out <= 16'h0383;    16'd25985: out <= 16'h0149;    16'd25986: out <= 16'h0670;    16'd25987: out <= 16'h0512;
    16'd25988: out <= 16'h0672;    16'd25989: out <= 16'h049E;    16'd25990: out <= 16'h088E;    16'd25991: out <= 16'h0162;
    16'd25992: out <= 16'h03AA;    16'd25993: out <= 16'h0587;    16'd25994: out <= 16'h07AA;    16'd25995: out <= 16'h0952;
    16'd25996: out <= 16'h0058;    16'd25997: out <= 16'h01DA;    16'd25998: out <= 16'h001F;    16'd25999: out <= 16'h00F7;
    16'd26000: out <= 16'h02BD;    16'd26001: out <= 16'h0625;    16'd26002: out <= 16'h0341;    16'd26003: out <= 16'hFDDC;
    16'd26004: out <= 16'h02D7;    16'd26005: out <= 16'h0407;    16'd26006: out <= 16'h029B;    16'd26007: out <= 16'h0A31;
    16'd26008: out <= 16'h049A;    16'd26009: out <= 16'h0101;    16'd26010: out <= 16'h0429;    16'd26011: out <= 16'h070E;
    16'd26012: out <= 16'h034D;    16'd26013: out <= 16'h0970;    16'd26014: out <= 16'hFA13;    16'd26015: out <= 16'hFE3E;
    16'd26016: out <= 16'h02C1;    16'd26017: out <= 16'h00B7;    16'd26018: out <= 16'hFCA9;    16'd26019: out <= 16'h0227;
    16'd26020: out <= 16'hFB7F;    16'd26021: out <= 16'h00C4;    16'd26022: out <= 16'h003C;    16'd26023: out <= 16'hFF05;
    16'd26024: out <= 16'hF573;    16'd26025: out <= 16'hFEB6;    16'd26026: out <= 16'h029A;    16'd26027: out <= 16'h00E8;
    16'd26028: out <= 16'h06E1;    16'd26029: out <= 16'hFA1C;    16'd26030: out <= 16'hFD9B;    16'd26031: out <= 16'h0232;
    16'd26032: out <= 16'hFB45;    16'd26033: out <= 16'h0234;    16'd26034: out <= 16'h00F7;    16'd26035: out <= 16'h051F;
    16'd26036: out <= 16'hFF9A;    16'd26037: out <= 16'hFFB2;    16'd26038: out <= 16'h0022;    16'd26039: out <= 16'hFEDF;
    16'd26040: out <= 16'h0517;    16'd26041: out <= 16'h02A8;    16'd26042: out <= 16'h09EE;    16'd26043: out <= 16'h0277;
    16'd26044: out <= 16'h0C0D;    16'd26045: out <= 16'h020C;    16'd26046: out <= 16'h099E;    16'd26047: out <= 16'h072D;
    16'd26048: out <= 16'h02A6;    16'd26049: out <= 16'h012F;    16'd26050: out <= 16'h02F8;    16'd26051: out <= 16'h07D9;
    16'd26052: out <= 16'hFE48;    16'd26053: out <= 16'hFBA4;    16'd26054: out <= 16'h055B;    16'd26055: out <= 16'h00B7;
    16'd26056: out <= 16'h0170;    16'd26057: out <= 16'h0501;    16'd26058: out <= 16'h0854;    16'd26059: out <= 16'h0672;
    16'd26060: out <= 16'h0BE6;    16'd26061: out <= 16'h08EF;    16'd26062: out <= 16'hFBF9;    16'd26063: out <= 16'h037E;
    16'd26064: out <= 16'h0783;    16'd26065: out <= 16'h0617;    16'd26066: out <= 16'h0798;    16'd26067: out <= 16'h0993;
    16'd26068: out <= 16'hFE9E;    16'd26069: out <= 16'h05CA;    16'd26070: out <= 16'h0817;    16'd26071: out <= 16'h0028;
    16'd26072: out <= 16'h060B;    16'd26073: out <= 16'hFCDA;    16'd26074: out <= 16'h0622;    16'd26075: out <= 16'h05E3;
    16'd26076: out <= 16'hF96A;    16'd26077: out <= 16'hFD25;    16'd26078: out <= 16'hFB26;    16'd26079: out <= 16'hFCDC;
    16'd26080: out <= 16'hF7D9;    16'd26081: out <= 16'h0330;    16'd26082: out <= 16'h035A;    16'd26083: out <= 16'h0020;
    16'd26084: out <= 16'hFC16;    16'd26085: out <= 16'hFA0E;    16'd26086: out <= 16'hF937;    16'd26087: out <= 16'h01EA;
    16'd26088: out <= 16'hF9A8;    16'd26089: out <= 16'hFE5B;    16'd26090: out <= 16'h0172;    16'd26091: out <= 16'hFBFE;
    16'd26092: out <= 16'hFC4A;    16'd26093: out <= 16'h0AD0;    16'd26094: out <= 16'hF840;    16'd26095: out <= 16'hFC73;
    16'd26096: out <= 16'hFDC4;    16'd26097: out <= 16'hFE13;    16'd26098: out <= 16'h025A;    16'd26099: out <= 16'h0172;
    16'd26100: out <= 16'h053B;    16'd26101: out <= 16'h018D;    16'd26102: out <= 16'hFEDD;    16'd26103: out <= 16'hFD12;
    16'd26104: out <= 16'hFE62;    16'd26105: out <= 16'h012A;    16'd26106: out <= 16'hF9C0;    16'd26107: out <= 16'h02F5;
    16'd26108: out <= 16'hFEA1;    16'd26109: out <= 16'hF848;    16'd26110: out <= 16'h00F7;    16'd26111: out <= 16'hFDE1;
    16'd26112: out <= 16'h0010;    16'd26113: out <= 16'hFF61;    16'd26114: out <= 16'hFEE9;    16'd26115: out <= 16'h07A7;
    16'd26116: out <= 16'hFC99;    16'd26117: out <= 16'h0151;    16'd26118: out <= 16'h0072;    16'd26119: out <= 16'h0072;
    16'd26120: out <= 16'hFB73;    16'd26121: out <= 16'h01D3;    16'd26122: out <= 16'hFD08;    16'd26123: out <= 16'hFD29;
    16'd26124: out <= 16'hFF98;    16'd26125: out <= 16'h00A0;    16'd26126: out <= 16'h0061;    16'd26127: out <= 16'hFB8F;
    16'd26128: out <= 16'hFF78;    16'd26129: out <= 16'hFEA1;    16'd26130: out <= 16'hFEC8;    16'd26131: out <= 16'h0259;
    16'd26132: out <= 16'hFF88;    16'd26133: out <= 16'hFFA5;    16'd26134: out <= 16'hFA4A;    16'd26135: out <= 16'hFCD0;
    16'd26136: out <= 16'h0870;    16'd26137: out <= 16'h05EB;    16'd26138: out <= 16'h017D;    16'd26139: out <= 16'h019B;
    16'd26140: out <= 16'h0412;    16'd26141: out <= 16'hFB53;    16'd26142: out <= 16'hFC53;    16'd26143: out <= 16'h08F7;
    16'd26144: out <= 16'h0486;    16'd26145: out <= 16'h081C;    16'd26146: out <= 16'h0209;    16'd26147: out <= 16'h07C3;
    16'd26148: out <= 16'hFF50;    16'd26149: out <= 16'h01DE;    16'd26150: out <= 16'h0373;    16'd26151: out <= 16'h03B0;
    16'd26152: out <= 16'hFF8F;    16'd26153: out <= 16'h0730;    16'd26154: out <= 16'h04DC;    16'd26155: out <= 16'h05B8;
    16'd26156: out <= 16'h071C;    16'd26157: out <= 16'hFEA6;    16'd26158: out <= 16'h0244;    16'd26159: out <= 16'h0340;
    16'd26160: out <= 16'h019E;    16'd26161: out <= 16'h025F;    16'd26162: out <= 16'h08FF;    16'd26163: out <= 16'h0252;
    16'd26164: out <= 16'h0199;    16'd26165: out <= 16'h050A;    16'd26166: out <= 16'h061A;    16'd26167: out <= 16'hFFAC;
    16'd26168: out <= 16'h07C5;    16'd26169: out <= 16'hFC8A;    16'd26170: out <= 16'h00ED;    16'd26171: out <= 16'h0AC1;
    16'd26172: out <= 16'h0AB4;    16'd26173: out <= 16'h05FE;    16'd26174: out <= 16'h054E;    16'd26175: out <= 16'h0025;
    16'd26176: out <= 16'h03D2;    16'd26177: out <= 16'h00E0;    16'd26178: out <= 16'h017C;    16'd26179: out <= 16'h0644;
    16'd26180: out <= 16'h0481;    16'd26181: out <= 16'h029D;    16'd26182: out <= 16'h0290;    16'd26183: out <= 16'h01AE;
    16'd26184: out <= 16'hFDC0;    16'd26185: out <= 16'h00F2;    16'd26186: out <= 16'hFEEE;    16'd26187: out <= 16'h0215;
    16'd26188: out <= 16'h0220;    16'd26189: out <= 16'hFD72;    16'd26190: out <= 16'hFF42;    16'd26191: out <= 16'h023B;
    16'd26192: out <= 16'hF847;    16'd26193: out <= 16'h0A24;    16'd26194: out <= 16'hFDA4;    16'd26195: out <= 16'h05CE;
    16'd26196: out <= 16'h0765;    16'd26197: out <= 16'hFECF;    16'd26198: out <= 16'hFE33;    16'd26199: out <= 16'h01F8;
    16'd26200: out <= 16'h08B1;    16'd26201: out <= 16'h0450;    16'd26202: out <= 16'h03BB;    16'd26203: out <= 16'h0299;
    16'd26204: out <= 16'h05BA;    16'd26205: out <= 16'h04F6;    16'd26206: out <= 16'hFFB6;    16'd26207: out <= 16'h0066;
    16'd26208: out <= 16'h03DD;    16'd26209: out <= 16'h0179;    16'd26210: out <= 16'h00DD;    16'd26211: out <= 16'hFC57;
    16'd26212: out <= 16'h0743;    16'd26213: out <= 16'h0490;    16'd26214: out <= 16'h0623;    16'd26215: out <= 16'hFBA5;
    16'd26216: out <= 16'h028F;    16'd26217: out <= 16'h0859;    16'd26218: out <= 16'h07B3;    16'd26219: out <= 16'h0394;
    16'd26220: out <= 16'h0480;    16'd26221: out <= 16'h07BA;    16'd26222: out <= 16'h0536;    16'd26223: out <= 16'h0371;
    16'd26224: out <= 16'hFE15;    16'd26225: out <= 16'hFE2C;    16'd26226: out <= 16'h08DE;    16'd26227: out <= 16'h0134;
    16'd26228: out <= 16'h0982;    16'd26229: out <= 16'h0C79;    16'd26230: out <= 16'h04D6;    16'd26231: out <= 16'h0652;
    16'd26232: out <= 16'h0273;    16'd26233: out <= 16'h022F;    16'd26234: out <= 16'hFF5A;    16'd26235: out <= 16'hFD7D;
    16'd26236: out <= 16'h00CB;    16'd26237: out <= 16'h00F4;    16'd26238: out <= 16'h0436;    16'd26239: out <= 16'hFEE6;
    16'd26240: out <= 16'h0836;    16'd26241: out <= 16'h0137;    16'd26242: out <= 16'h03D4;    16'd26243: out <= 16'h056F;
    16'd26244: out <= 16'h0192;    16'd26245: out <= 16'h0583;    16'd26246: out <= 16'hFC43;    16'd26247: out <= 16'h04AD;
    16'd26248: out <= 16'h0676;    16'd26249: out <= 16'h079E;    16'd26250: out <= 16'h045F;    16'd26251: out <= 16'hFB49;
    16'd26252: out <= 16'h0440;    16'd26253: out <= 16'h0132;    16'd26254: out <= 16'h06A9;    16'd26255: out <= 16'h0766;
    16'd26256: out <= 16'h077E;    16'd26257: out <= 16'h042B;    16'd26258: out <= 16'h07B4;    16'd26259: out <= 16'hFB7A;
    16'd26260: out <= 16'hFF1B;    16'd26261: out <= 16'hFFD4;    16'd26262: out <= 16'h0957;    16'd26263: out <= 16'h032C;
    16'd26264: out <= 16'h04F3;    16'd26265: out <= 16'h058C;    16'd26266: out <= 16'h03E6;    16'd26267: out <= 16'h02A9;
    16'd26268: out <= 16'h084A;    16'd26269: out <= 16'h01F4;    16'd26270: out <= 16'h0B99;    16'd26271: out <= 16'hFD92;
    16'd26272: out <= 16'hFFB2;    16'd26273: out <= 16'h056F;    16'd26274: out <= 16'h04E7;    16'd26275: out <= 16'hFEB3;
    16'd26276: out <= 16'hFE58;    16'd26277: out <= 16'h0015;    16'd26278: out <= 16'hF8FA;    16'd26279: out <= 16'h0078;
    16'd26280: out <= 16'hFDB4;    16'd26281: out <= 16'hF7C4;    16'd26282: out <= 16'hFEEE;    16'd26283: out <= 16'h00C4;
    16'd26284: out <= 16'h0499;    16'd26285: out <= 16'hFC77;    16'd26286: out <= 16'hFAEB;    16'd26287: out <= 16'h0507;
    16'd26288: out <= 16'h00DC;    16'd26289: out <= 16'h02A4;    16'd26290: out <= 16'h069E;    16'd26291: out <= 16'h095C;
    16'd26292: out <= 16'h08CD;    16'd26293: out <= 16'h081E;    16'd26294: out <= 16'h018E;    16'd26295: out <= 16'h08AE;
    16'd26296: out <= 16'h01F0;    16'd26297: out <= 16'h021F;    16'd26298: out <= 16'h097D;    16'd26299: out <= 16'h0175;
    16'd26300: out <= 16'h0A20;    16'd26301: out <= 16'h0033;    16'd26302: out <= 16'h031B;    16'd26303: out <= 16'h03D4;
    16'd26304: out <= 16'h041D;    16'd26305: out <= 16'h0272;    16'd26306: out <= 16'h0BD1;    16'd26307: out <= 16'h03CF;
    16'd26308: out <= 16'hFC8F;    16'd26309: out <= 16'h0181;    16'd26310: out <= 16'h0660;    16'd26311: out <= 16'h0913;
    16'd26312: out <= 16'hFF1A;    16'd26313: out <= 16'h00D4;    16'd26314: out <= 16'h0035;    16'd26315: out <= 16'hFE82;
    16'd26316: out <= 16'h0205;    16'd26317: out <= 16'h03AE;    16'd26318: out <= 16'h074B;    16'd26319: out <= 16'h0868;
    16'd26320: out <= 16'h0B17;    16'd26321: out <= 16'h029F;    16'd26322: out <= 16'h08CA;    16'd26323: out <= 16'h0310;
    16'd26324: out <= 16'hFD35;    16'd26325: out <= 16'h0763;    16'd26326: out <= 16'hFDBC;    16'd26327: out <= 16'h0369;
    16'd26328: out <= 16'h054A;    16'd26329: out <= 16'h0619;    16'd26330: out <= 16'h02C5;    16'd26331: out <= 16'h0205;
    16'd26332: out <= 16'hFD32;    16'd26333: out <= 16'hFF2F;    16'd26334: out <= 16'h05C4;    16'd26335: out <= 16'hFFB0;
    16'd26336: out <= 16'hF98A;    16'd26337: out <= 16'h0211;    16'd26338: out <= 16'h039D;    16'd26339: out <= 16'hFD0A;
    16'd26340: out <= 16'hFC8B;    16'd26341: out <= 16'h0731;    16'd26342: out <= 16'hFBE0;    16'd26343: out <= 16'h0637;
    16'd26344: out <= 16'h06EA;    16'd26345: out <= 16'h0289;    16'd26346: out <= 16'hFEC3;    16'd26347: out <= 16'h019B;
    16'd26348: out <= 16'h0187;    16'd26349: out <= 16'hFDBE;    16'd26350: out <= 16'hFF01;    16'd26351: out <= 16'h0668;
    16'd26352: out <= 16'hFD45;    16'd26353: out <= 16'hFE5E;    16'd26354: out <= 16'h0408;    16'd26355: out <= 16'hFF4B;
    16'd26356: out <= 16'hFE0F;    16'd26357: out <= 16'h06D2;    16'd26358: out <= 16'h00D1;    16'd26359: out <= 16'hFD97;
    16'd26360: out <= 16'h0133;    16'd26361: out <= 16'h0461;    16'd26362: out <= 16'hFDD0;    16'd26363: out <= 16'hFE93;
    16'd26364: out <= 16'hFEBA;    16'd26365: out <= 16'h0112;    16'd26366: out <= 16'hFDF4;    16'd26367: out <= 16'hFCC0;
    16'd26368: out <= 16'hFE66;    16'd26369: out <= 16'h00B7;    16'd26370: out <= 16'hFCC7;    16'd26371: out <= 16'h0068;
    16'd26372: out <= 16'hF8DE;    16'd26373: out <= 16'hFD69;    16'd26374: out <= 16'h0148;    16'd26375: out <= 16'hFE8B;
    16'd26376: out <= 16'h00AC;    16'd26377: out <= 16'h06BF;    16'd26378: out <= 16'hFBE9;    16'd26379: out <= 16'h0055;
    16'd26380: out <= 16'hFE75;    16'd26381: out <= 16'h0234;    16'd26382: out <= 16'hFDDB;    16'd26383: out <= 16'h035D;
    16'd26384: out <= 16'h009D;    16'd26385: out <= 16'h052B;    16'd26386: out <= 16'hFE6C;    16'd26387: out <= 16'h059B;
    16'd26388: out <= 16'hFCFB;    16'd26389: out <= 16'hFE1A;    16'd26390: out <= 16'h07C5;    16'd26391: out <= 16'h047F;
    16'd26392: out <= 16'hFFC0;    16'd26393: out <= 16'h0135;    16'd26394: out <= 16'hFEE3;    16'd26395: out <= 16'h0160;
    16'd26396: out <= 16'hFEBE;    16'd26397: out <= 16'hFAB6;    16'd26398: out <= 16'hFF0F;    16'd26399: out <= 16'h06A4;
    16'd26400: out <= 16'h032F;    16'd26401: out <= 16'h048D;    16'd26402: out <= 16'h058E;    16'd26403: out <= 16'h01EA;
    16'd26404: out <= 16'h04F1;    16'd26405: out <= 16'h03E0;    16'd26406: out <= 16'h09BA;    16'd26407: out <= 16'h009B;
    16'd26408: out <= 16'h0379;    16'd26409: out <= 16'h0031;    16'd26410: out <= 16'h05E7;    16'd26411: out <= 16'h0869;
    16'd26412: out <= 16'hFE12;    16'd26413: out <= 16'h03BB;    16'd26414: out <= 16'h05EA;    16'd26415: out <= 16'h0856;
    16'd26416: out <= 16'h0461;    16'd26417: out <= 16'h08DD;    16'd26418: out <= 16'h0707;    16'd26419: out <= 16'h01D9;
    16'd26420: out <= 16'h0042;    16'd26421: out <= 16'h0068;    16'd26422: out <= 16'h0637;    16'd26423: out <= 16'h0641;
    16'd26424: out <= 16'h020B;    16'd26425: out <= 16'h00B9;    16'd26426: out <= 16'h02CC;    16'd26427: out <= 16'hFD94;
    16'd26428: out <= 16'hFC31;    16'd26429: out <= 16'h0462;    16'd26430: out <= 16'h09BA;    16'd26431: out <= 16'h050C;
    16'd26432: out <= 16'h0286;    16'd26433: out <= 16'h001D;    16'd26434: out <= 16'h03B4;    16'd26435: out <= 16'hFADE;
    16'd26436: out <= 16'h07E9;    16'd26437: out <= 16'h052E;    16'd26438: out <= 16'h0959;    16'd26439: out <= 16'h00D8;
    16'd26440: out <= 16'hFE56;    16'd26441: out <= 16'hFC94;    16'd26442: out <= 16'hFF9F;    16'd26443: out <= 16'h04D3;
    16'd26444: out <= 16'hFF82;    16'd26445: out <= 16'h0563;    16'd26446: out <= 16'hFCD4;    16'd26447: out <= 16'h04BD;
    16'd26448: out <= 16'h0163;    16'd26449: out <= 16'h03FF;    16'd26450: out <= 16'h011B;    16'd26451: out <= 16'h05E8;
    16'd26452: out <= 16'h08CE;    16'd26453: out <= 16'hFC21;    16'd26454: out <= 16'h060F;    16'd26455: out <= 16'h030D;
    16'd26456: out <= 16'hFC30;    16'd26457: out <= 16'h02DB;    16'd26458: out <= 16'h05D1;    16'd26459: out <= 16'h005B;
    16'd26460: out <= 16'hFC09;    16'd26461: out <= 16'h0439;    16'd26462: out <= 16'h076B;    16'd26463: out <= 16'h0640;
    16'd26464: out <= 16'h0715;    16'd26465: out <= 16'hFED3;    16'd26466: out <= 16'h0670;    16'd26467: out <= 16'h004C;
    16'd26468: out <= 16'h0374;    16'd26469: out <= 16'h003D;    16'd26470: out <= 16'hFF81;    16'd26471: out <= 16'h071C;
    16'd26472: out <= 16'h0357;    16'd26473: out <= 16'h049E;    16'd26474: out <= 16'hFE21;    16'd26475: out <= 16'h0919;
    16'd26476: out <= 16'h0684;    16'd26477: out <= 16'h02B3;    16'd26478: out <= 16'h08BD;    16'd26479: out <= 16'hFFC6;
    16'd26480: out <= 16'h02C4;    16'd26481: out <= 16'h022E;    16'd26482: out <= 16'h07D2;    16'd26483: out <= 16'h0A23;
    16'd26484: out <= 16'h092E;    16'd26485: out <= 16'h02B8;    16'd26486: out <= 16'h0124;    16'd26487: out <= 16'h0724;
    16'd26488: out <= 16'h0453;    16'd26489: out <= 16'h0510;    16'd26490: out <= 16'h014F;    16'd26491: out <= 16'h0BA6;
    16'd26492: out <= 16'h0119;    16'd26493: out <= 16'h065D;    16'd26494: out <= 16'hFEE7;    16'd26495: out <= 16'h00D7;
    16'd26496: out <= 16'h0C1A;    16'd26497: out <= 16'hFE83;    16'd26498: out <= 16'h04E3;    16'd26499: out <= 16'h076E;
    16'd26500: out <= 16'hFF31;    16'd26501: out <= 16'h023A;    16'd26502: out <= 16'hFD50;    16'd26503: out <= 16'h015E;
    16'd26504: out <= 16'hFCD9;    16'd26505: out <= 16'h0497;    16'd26506: out <= 16'h07A3;    16'd26507: out <= 16'h04A9;
    16'd26508: out <= 16'h05B9;    16'd26509: out <= 16'h0360;    16'd26510: out <= 16'h0549;    16'd26511: out <= 16'h0644;
    16'd26512: out <= 16'h01DA;    16'd26513: out <= 16'hFDDA;    16'd26514: out <= 16'h033D;    16'd26515: out <= 16'h05FB;
    16'd26516: out <= 16'h05D5;    16'd26517: out <= 16'hFCFE;    16'd26518: out <= 16'h0865;    16'd26519: out <= 16'hFA29;
    16'd26520: out <= 16'h04DC;    16'd26521: out <= 16'h0031;    16'd26522: out <= 16'h04E0;    16'd26523: out <= 16'h05B2;
    16'd26524: out <= 16'h0488;    16'd26525: out <= 16'h0F44;    16'd26526: out <= 16'h0278;    16'd26527: out <= 16'hFEBF;
    16'd26528: out <= 16'h069E;    16'd26529: out <= 16'h015C;    16'd26530: out <= 16'hFF9B;    16'd26531: out <= 16'hFE0E;
    16'd26532: out <= 16'hFD80;    16'd26533: out <= 16'h00E5;    16'd26534: out <= 16'hFEAA;    16'd26535: out <= 16'hF836;
    16'd26536: out <= 16'hFF1B;    16'd26537: out <= 16'h017C;    16'd26538: out <= 16'h035E;    16'd26539: out <= 16'h04CF;
    16'd26540: out <= 16'h002B;    16'd26541: out <= 16'hFE08;    16'd26542: out <= 16'h0110;    16'd26543: out <= 16'h01CB;
    16'd26544: out <= 16'h0625;    16'd26545: out <= 16'hFF47;    16'd26546: out <= 16'h086A;    16'd26547: out <= 16'hFD93;
    16'd26548: out <= 16'hFBB3;    16'd26549: out <= 16'hFDE6;    16'd26550: out <= 16'h0530;    16'd26551: out <= 16'hFF26;
    16'd26552: out <= 16'h006B;    16'd26553: out <= 16'h023C;    16'd26554: out <= 16'h0510;    16'd26555: out <= 16'h0136;
    16'd26556: out <= 16'hFDD7;    16'd26557: out <= 16'h04D9;    16'd26558: out <= 16'hFCA1;    16'd26559: out <= 16'h0480;
    16'd26560: out <= 16'h0266;    16'd26561: out <= 16'hFC53;    16'd26562: out <= 16'h06CD;    16'd26563: out <= 16'h018F;
    16'd26564: out <= 16'h02E4;    16'd26565: out <= 16'h08B8;    16'd26566: out <= 16'h0563;    16'd26567: out <= 16'h0693;
    16'd26568: out <= 16'h0369;    16'd26569: out <= 16'h067C;    16'd26570: out <= 16'h007B;    16'd26571: out <= 16'hF9F2;
    16'd26572: out <= 16'h0E70;    16'd26573: out <= 16'h06C7;    16'd26574: out <= 16'h0752;    16'd26575: out <= 16'h062B;
    16'd26576: out <= 16'h0518;    16'd26577: out <= 16'h037E;    16'd26578: out <= 16'hFF10;    16'd26579: out <= 16'h0B38;
    16'd26580: out <= 16'h0451;    16'd26581: out <= 16'h0A25;    16'd26582: out <= 16'h0293;    16'd26583: out <= 16'h06E1;
    16'd26584: out <= 16'h0230;    16'd26585: out <= 16'h0115;    16'd26586: out <= 16'hFC28;    16'd26587: out <= 16'h0552;
    16'd26588: out <= 16'hF943;    16'd26589: out <= 16'hFE7B;    16'd26590: out <= 16'hF980;    16'd26591: out <= 16'h07B4;
    16'd26592: out <= 16'hFD3D;    16'd26593: out <= 16'hFE41;    16'd26594: out <= 16'h00C8;    16'd26595: out <= 16'h0761;
    16'd26596: out <= 16'hFCB2;    16'd26597: out <= 16'hF9EF;    16'd26598: out <= 16'h03AA;    16'd26599: out <= 16'h0031;
    16'd26600: out <= 16'h0066;    16'd26601: out <= 16'h0243;    16'd26602: out <= 16'hFE42;    16'd26603: out <= 16'hFF13;
    16'd26604: out <= 16'hFF95;    16'd26605: out <= 16'h023C;    16'd26606: out <= 16'hF9AB;    16'd26607: out <= 16'hF9D8;
    16'd26608: out <= 16'hF895;    16'd26609: out <= 16'h0056;    16'd26610: out <= 16'h04DC;    16'd26611: out <= 16'hFA25;
    16'd26612: out <= 16'hFFBC;    16'd26613: out <= 16'hFCE6;    16'd26614: out <= 16'h062D;    16'd26615: out <= 16'hFF69;
    16'd26616: out <= 16'hFC85;    16'd26617: out <= 16'h022C;    16'd26618: out <= 16'h06DE;    16'd26619: out <= 16'h03CE;
    16'd26620: out <= 16'h0027;    16'd26621: out <= 16'h0803;    16'd26622: out <= 16'h0168;    16'd26623: out <= 16'hFE8F;
    16'd26624: out <= 16'hFD76;    16'd26625: out <= 16'h0564;    16'd26626: out <= 16'hFCF5;    16'd26627: out <= 16'h041A;
    16'd26628: out <= 16'hFA14;    16'd26629: out <= 16'hFFC3;    16'd26630: out <= 16'h031B;    16'd26631: out <= 16'hFF52;
    16'd26632: out <= 16'h0183;    16'd26633: out <= 16'h00DD;    16'd26634: out <= 16'hFDFD;    16'd26635: out <= 16'h028C;
    16'd26636: out <= 16'hFB70;    16'd26637: out <= 16'hFBF7;    16'd26638: out <= 16'h02C5;    16'd26639: out <= 16'h00B5;
    16'd26640: out <= 16'h0299;    16'd26641: out <= 16'hF5AD;    16'd26642: out <= 16'hF8E2;    16'd26643: out <= 16'hFD94;
    16'd26644: out <= 16'hFDB0;    16'd26645: out <= 16'hFFA8;    16'd26646: out <= 16'h03A8;    16'd26647: out <= 16'hFFC5;
    16'd26648: out <= 16'hF8AE;    16'd26649: out <= 16'h0020;    16'd26650: out <= 16'h02A7;    16'd26651: out <= 16'h064F;
    16'd26652: out <= 16'h03A7;    16'd26653: out <= 16'hFD40;    16'd26654: out <= 16'hFE85;    16'd26655: out <= 16'h02E4;
    16'd26656: out <= 16'h0A12;    16'd26657: out <= 16'h0A6F;    16'd26658: out <= 16'h0000;    16'd26659: out <= 16'h041F;
    16'd26660: out <= 16'h0274;    16'd26661: out <= 16'h038C;    16'd26662: out <= 16'h04DB;    16'd26663: out <= 16'h08EF;
    16'd26664: out <= 16'h03F5;    16'd26665: out <= 16'hFE53;    16'd26666: out <= 16'h0551;    16'd26667: out <= 16'h0D34;
    16'd26668: out <= 16'h06FC;    16'd26669: out <= 16'hFFBF;    16'd26670: out <= 16'h03A6;    16'd26671: out <= 16'h04CF;
    16'd26672: out <= 16'h0339;    16'd26673: out <= 16'h019A;    16'd26674: out <= 16'h0422;    16'd26675: out <= 16'h0389;
    16'd26676: out <= 16'h0484;    16'd26677: out <= 16'h048F;    16'd26678: out <= 16'h043B;    16'd26679: out <= 16'h00BC;
    16'd26680: out <= 16'h0174;    16'd26681: out <= 16'h065E;    16'd26682: out <= 16'h012D;    16'd26683: out <= 16'h0024;
    16'd26684: out <= 16'h033B;    16'd26685: out <= 16'hFA51;    16'd26686: out <= 16'h016E;    16'd26687: out <= 16'h0534;
    16'd26688: out <= 16'h01EC;    16'd26689: out <= 16'h05AA;    16'd26690: out <= 16'h0887;    16'd26691: out <= 16'h064A;
    16'd26692: out <= 16'h04E0;    16'd26693: out <= 16'h0869;    16'd26694: out <= 16'h06A2;    16'd26695: out <= 16'h002C;
    16'd26696: out <= 16'h00D5;    16'd26697: out <= 16'h0300;    16'd26698: out <= 16'h0300;    16'd26699: out <= 16'hFD46;
    16'd26700: out <= 16'h0271;    16'd26701: out <= 16'h033B;    16'd26702: out <= 16'h045F;    16'd26703: out <= 16'h00D0;
    16'd26704: out <= 16'h00E2;    16'd26705: out <= 16'h0AFA;    16'd26706: out <= 16'h0525;    16'd26707: out <= 16'hFED3;
    16'd26708: out <= 16'h0336;    16'd26709: out <= 16'h056E;    16'd26710: out <= 16'h0673;    16'd26711: out <= 16'h03D9;
    16'd26712: out <= 16'h077E;    16'd26713: out <= 16'h035A;    16'd26714: out <= 16'h01C0;    16'd26715: out <= 16'h07E4;
    16'd26716: out <= 16'h07B6;    16'd26717: out <= 16'h04D7;    16'd26718: out <= 16'h03C7;    16'd26719: out <= 16'h03C3;
    16'd26720: out <= 16'h0546;    16'd26721: out <= 16'h0469;    16'd26722: out <= 16'h038E;    16'd26723: out <= 16'h01F2;
    16'd26724: out <= 16'h013F;    16'd26725: out <= 16'h07F6;    16'd26726: out <= 16'h0606;    16'd26727: out <= 16'h04E4;
    16'd26728: out <= 16'hFBCD;    16'd26729: out <= 16'hFD59;    16'd26730: out <= 16'h0091;    16'd26731: out <= 16'h05C3;
    16'd26732: out <= 16'h022F;    16'd26733: out <= 16'h02B6;    16'd26734: out <= 16'h059B;    16'd26735: out <= 16'hFDF5;
    16'd26736: out <= 16'h0377;    16'd26737: out <= 16'hFDF7;    16'd26738: out <= 16'h073C;    16'd26739: out <= 16'h0603;
    16'd26740: out <= 16'h02DD;    16'd26741: out <= 16'h07D0;    16'd26742: out <= 16'h09BE;    16'd26743: out <= 16'h0200;
    16'd26744: out <= 16'hFD97;    16'd26745: out <= 16'h00F8;    16'd26746: out <= 16'h01E1;    16'd26747: out <= 16'h0A6A;
    16'd26748: out <= 16'h0A8D;    16'd26749: out <= 16'h0930;    16'd26750: out <= 16'h07DA;    16'd26751: out <= 16'hFFF0;
    16'd26752: out <= 16'h024E;    16'd26753: out <= 16'h0446;    16'd26754: out <= 16'h0355;    16'd26755: out <= 16'hFEB6;
    16'd26756: out <= 16'h034E;    16'd26757: out <= 16'h004C;    16'd26758: out <= 16'h01C7;    16'd26759: out <= 16'h00E1;
    16'd26760: out <= 16'h02C8;    16'd26761: out <= 16'h01C1;    16'd26762: out <= 16'h0975;    16'd26763: out <= 16'h01A6;
    16'd26764: out <= 16'h02A2;    16'd26765: out <= 16'h0484;    16'd26766: out <= 16'h00D9;    16'd26767: out <= 16'h0421;
    16'd26768: out <= 16'h07B2;    16'd26769: out <= 16'h07B0;    16'd26770: out <= 16'h02E1;    16'd26771: out <= 16'h045B;
    16'd26772: out <= 16'h02C1;    16'd26773: out <= 16'h08EC;    16'd26774: out <= 16'h015A;    16'd26775: out <= 16'h064A;
    16'd26776: out <= 16'hFFD4;    16'd26777: out <= 16'hFBF3;    16'd26778: out <= 16'h0079;    16'd26779: out <= 16'h0825;
    16'd26780: out <= 16'h05E2;    16'd26781: out <= 16'h076B;    16'd26782: out <= 16'h01DC;    16'd26783: out <= 16'h04B1;
    16'd26784: out <= 16'h080C;    16'd26785: out <= 16'hFE50;    16'd26786: out <= 16'h0283;    16'd26787: out <= 16'h03A0;
    16'd26788: out <= 16'hFC13;    16'd26789: out <= 16'hFF63;    16'd26790: out <= 16'h0644;    16'd26791: out <= 16'hF854;
    16'd26792: out <= 16'h012F;    16'd26793: out <= 16'h020F;    16'd26794: out <= 16'hFC31;    16'd26795: out <= 16'hFE3B;
    16'd26796: out <= 16'hFC94;    16'd26797: out <= 16'h0415;    16'd26798: out <= 16'hFD94;    16'd26799: out <= 16'hFB0A;
    16'd26800: out <= 16'h01F8;    16'd26801: out <= 16'hF962;    16'd26802: out <= 16'hFC0D;    16'd26803: out <= 16'hFF8B;
    16'd26804: out <= 16'h04E5;    16'd26805: out <= 16'h0C6C;    16'd26806: out <= 16'hFB45;    16'd26807: out <= 16'hFF61;
    16'd26808: out <= 16'h075C;    16'd26809: out <= 16'h0333;    16'd26810: out <= 16'h002B;    16'd26811: out <= 16'h02D2;
    16'd26812: out <= 16'hFFEB;    16'd26813: out <= 16'h0496;    16'd26814: out <= 16'hFC5D;    16'd26815: out <= 16'hFF4A;
    16'd26816: out <= 16'h0190;    16'd26817: out <= 16'h04A5;    16'd26818: out <= 16'h018C;    16'd26819: out <= 16'h023F;
    16'd26820: out <= 16'h01EC;    16'd26821: out <= 16'h0042;    16'd26822: out <= 16'hFA96;    16'd26823: out <= 16'h071E;
    16'd26824: out <= 16'h0280;    16'd26825: out <= 16'h089B;    16'd26826: out <= 16'h04B5;    16'd26827: out <= 16'h0BBB;
    16'd26828: out <= 16'h03C3;    16'd26829: out <= 16'hFEEB;    16'd26830: out <= 16'h0955;    16'd26831: out <= 16'h04F8;
    16'd26832: out <= 16'h0805;    16'd26833: out <= 16'h07F6;    16'd26834: out <= 16'h0351;    16'd26835: out <= 16'h02FA;
    16'd26836: out <= 16'h0591;    16'd26837: out <= 16'h02F4;    16'd26838: out <= 16'h0356;    16'd26839: out <= 16'h091A;
    16'd26840: out <= 16'h0253;    16'd26841: out <= 16'hFE3A;    16'd26842: out <= 16'h0539;    16'd26843: out <= 16'hFE87;
    16'd26844: out <= 16'h0187;    16'd26845: out <= 16'h0013;    16'd26846: out <= 16'h01A9;    16'd26847: out <= 16'h0331;
    16'd26848: out <= 16'h006B;    16'd26849: out <= 16'hFF03;    16'd26850: out <= 16'hFB4F;    16'd26851: out <= 16'hF78C;
    16'd26852: out <= 16'hFFAB;    16'd26853: out <= 16'h0795;    16'd26854: out <= 16'hFF89;    16'd26855: out <= 16'hFF4A;
    16'd26856: out <= 16'h0154;    16'd26857: out <= 16'hFE0F;    16'd26858: out <= 16'hF6D7;    16'd26859: out <= 16'hFBC3;
    16'd26860: out <= 16'h046D;    16'd26861: out <= 16'h0293;    16'd26862: out <= 16'hFBC2;    16'd26863: out <= 16'hF988;
    16'd26864: out <= 16'hFE1E;    16'd26865: out <= 16'h010A;    16'd26866: out <= 16'h04A5;    16'd26867: out <= 16'h0286;
    16'd26868: out <= 16'h0130;    16'd26869: out <= 16'h0038;    16'd26870: out <= 16'hFFD1;    16'd26871: out <= 16'h0219;
    16'd26872: out <= 16'hFE8B;    16'd26873: out <= 16'hFE84;    16'd26874: out <= 16'h0296;    16'd26875: out <= 16'h016A;
    16'd26876: out <= 16'h045F;    16'd26877: out <= 16'h00C4;    16'd26878: out <= 16'hFE99;    16'd26879: out <= 16'hFF7A;
    16'd26880: out <= 16'hFFCA;    16'd26881: out <= 16'hFC98;    16'd26882: out <= 16'h018F;    16'd26883: out <= 16'h08DF;
    16'd26884: out <= 16'h00B7;    16'd26885: out <= 16'h05DD;    16'd26886: out <= 16'hFE59;    16'd26887: out <= 16'hF9C9;
    16'd26888: out <= 16'hFE3D;    16'd26889: out <= 16'h0352;    16'd26890: out <= 16'hF841;    16'd26891: out <= 16'h0290;
    16'd26892: out <= 16'h014F;    16'd26893: out <= 16'h045D;    16'd26894: out <= 16'h00A0;    16'd26895: out <= 16'hFD22;
    16'd26896: out <= 16'hFC91;    16'd26897: out <= 16'hFCAF;    16'd26898: out <= 16'hF90F;    16'd26899: out <= 16'hFEBB;
    16'd26900: out <= 16'hFEF6;    16'd26901: out <= 16'hFECC;    16'd26902: out <= 16'hFD79;    16'd26903: out <= 16'h01C0;
    16'd26904: out <= 16'h015B;    16'd26905: out <= 16'h072E;    16'd26906: out <= 16'hFAB1;    16'd26907: out <= 16'hFB88;
    16'd26908: out <= 16'h03F1;    16'd26909: out <= 16'h021D;    16'd26910: out <= 16'hFC55;    16'd26911: out <= 16'hF8F3;
    16'd26912: out <= 16'h0419;    16'd26913: out <= 16'h082B;    16'd26914: out <= 16'h0608;    16'd26915: out <= 16'h08B1;
    16'd26916: out <= 16'h0442;    16'd26917: out <= 16'h07DE;    16'd26918: out <= 16'h045B;    16'd26919: out <= 16'h06A7;
    16'd26920: out <= 16'hFD26;    16'd26921: out <= 16'h0584;    16'd26922: out <= 16'h02F0;    16'd26923: out <= 16'hFE58;
    16'd26924: out <= 16'h03B0;    16'd26925: out <= 16'h0864;    16'd26926: out <= 16'hFE46;    16'd26927: out <= 16'h0420;
    16'd26928: out <= 16'h0505;    16'd26929: out <= 16'h01F7;    16'd26930: out <= 16'h0214;    16'd26931: out <= 16'h05D3;
    16'd26932: out <= 16'h0186;    16'd26933: out <= 16'h0010;    16'd26934: out <= 16'h094A;    16'd26935: out <= 16'h0531;
    16'd26936: out <= 16'h0206;    16'd26937: out <= 16'h05DD;    16'd26938: out <= 16'h0803;    16'd26939: out <= 16'h08C0;
    16'd26940: out <= 16'hFFD2;    16'd26941: out <= 16'h0268;    16'd26942: out <= 16'h0083;    16'd26943: out <= 16'h02CA;
    16'd26944: out <= 16'h012A;    16'd26945: out <= 16'h05A5;    16'd26946: out <= 16'h03D7;    16'd26947: out <= 16'h03BF;
    16'd26948: out <= 16'hFEE6;    16'd26949: out <= 16'h0594;    16'd26950: out <= 16'h08FA;    16'd26951: out <= 16'h0799;
    16'd26952: out <= 16'hFDC8;    16'd26953: out <= 16'h06F3;    16'd26954: out <= 16'h01D9;    16'd26955: out <= 16'h06CF;
    16'd26956: out <= 16'hF752;    16'd26957: out <= 16'h094B;    16'd26958: out <= 16'h05CA;    16'd26959: out <= 16'h05DD;
    16'd26960: out <= 16'h08B8;    16'd26961: out <= 16'h020E;    16'd26962: out <= 16'h042F;    16'd26963: out <= 16'h0149;
    16'd26964: out <= 16'h08A1;    16'd26965: out <= 16'hFEA6;    16'd26966: out <= 16'h0B24;    16'd26967: out <= 16'hFE64;
    16'd26968: out <= 16'h0287;    16'd26969: out <= 16'h01A0;    16'd26970: out <= 16'h03AF;    16'd26971: out <= 16'h03BB;
    16'd26972: out <= 16'h0D2D;    16'd26973: out <= 16'h00D0;    16'd26974: out <= 16'h035A;    16'd26975: out <= 16'h05B6;
    16'd26976: out <= 16'h0901;    16'd26977: out <= 16'h065A;    16'd26978: out <= 16'h024C;    16'd26979: out <= 16'hFF32;
    16'd26980: out <= 16'hFCB7;    16'd26981: out <= 16'h08DF;    16'd26982: out <= 16'h00ED;    16'd26983: out <= 16'h0135;
    16'd26984: out <= 16'h01C4;    16'd26985: out <= 16'h00B6;    16'd26986: out <= 16'h06AB;    16'd26987: out <= 16'h062A;
    16'd26988: out <= 16'h01A5;    16'd26989: out <= 16'h04B4;    16'd26990: out <= 16'hFCCB;    16'd26991: out <= 16'hFEF5;
    16'd26992: out <= 16'h0102;    16'd26993: out <= 16'h01F0;    16'd26994: out <= 16'h0404;    16'd26995: out <= 16'h0777;
    16'd26996: out <= 16'h0487;    16'd26997: out <= 16'h0734;    16'd26998: out <= 16'h0334;    16'd26999: out <= 16'h03D5;
    16'd27000: out <= 16'hFFB0;    16'd27001: out <= 16'h0442;    16'd27002: out <= 16'h07D5;    16'd27003: out <= 16'h0424;
    16'd27004: out <= 16'h0812;    16'd27005: out <= 16'h056F;    16'd27006: out <= 16'h06F9;    16'd27007: out <= 16'h0878;
    16'd27008: out <= 16'hFFE2;    16'd27009: out <= 16'h04AB;    16'd27010: out <= 16'h035B;    16'd27011: out <= 16'h02E6;
    16'd27012: out <= 16'h0440;    16'd27013: out <= 16'h061A;    16'd27014: out <= 16'h03B2;    16'd27015: out <= 16'h0669;
    16'd27016: out <= 16'h0515;    16'd27017: out <= 16'h04DA;    16'd27018: out <= 16'hFF4A;    16'd27019: out <= 16'h0041;
    16'd27020: out <= 16'h0A87;    16'd27021: out <= 16'h054F;    16'd27022: out <= 16'h0510;    16'd27023: out <= 16'h0996;
    16'd27024: out <= 16'hFDD7;    16'd27025: out <= 16'h07BE;    16'd27026: out <= 16'h0727;    16'd27027: out <= 16'h0109;
    16'd27028: out <= 16'h0129;    16'd27029: out <= 16'h0608;    16'd27030: out <= 16'h004D;    16'd27031: out <= 16'h047A;
    16'd27032: out <= 16'h011D;    16'd27033: out <= 16'h06C0;    16'd27034: out <= 16'h05D9;    16'd27035: out <= 16'h0800;
    16'd27036: out <= 16'hFC72;    16'd27037: out <= 16'h0009;    16'd27038: out <= 16'h0750;    16'd27039: out <= 16'hFFFA;
    16'd27040: out <= 16'h03BF;    16'd27041: out <= 16'h056E;    16'd27042: out <= 16'h074C;    16'd27043: out <= 16'hFA2E;
    16'd27044: out <= 16'hF8D5;    16'd27045: out <= 16'hFBC0;    16'd27046: out <= 16'hFEE3;    16'd27047: out <= 16'hFC22;
    16'd27048: out <= 16'h0136;    16'd27049: out <= 16'hFAAC;    16'd27050: out <= 16'h01A9;    16'd27051: out <= 16'hF916;
    16'd27052: out <= 16'h04C4;    16'd27053: out <= 16'h02E1;    16'd27054: out <= 16'hFE36;    16'd27055: out <= 16'hF91A;
    16'd27056: out <= 16'h06C4;    16'd27057: out <= 16'h06F2;    16'd27058: out <= 16'h0217;    16'd27059: out <= 16'hFF79;
    16'd27060: out <= 16'h04EB;    16'd27061: out <= 16'h0033;    16'd27062: out <= 16'h0173;    16'd27063: out <= 16'h0041;
    16'd27064: out <= 16'hFE26;    16'd27065: out <= 16'h069B;    16'd27066: out <= 16'h01F5;    16'd27067: out <= 16'h0CFD;
    16'd27068: out <= 16'hFF6A;    16'd27069: out <= 16'h05FA;    16'd27070: out <= 16'h07B8;    16'd27071: out <= 16'h043A;
    16'd27072: out <= 16'h04FA;    16'd27073: out <= 16'h02CA;    16'd27074: out <= 16'h04A4;    16'd27075: out <= 16'h0305;
    16'd27076: out <= 16'h053F;    16'd27077: out <= 16'h0847;    16'd27078: out <= 16'hFF94;    16'd27079: out <= 16'h0601;
    16'd27080: out <= 16'h0320;    16'd27081: out <= 16'hFF1E;    16'd27082: out <= 16'h01C8;    16'd27083: out <= 16'h0441;
    16'd27084: out <= 16'h0188;    16'd27085: out <= 16'h0062;    16'd27086: out <= 16'h0182;    16'd27087: out <= 16'h02EA;
    16'd27088: out <= 16'h07A0;    16'd27089: out <= 16'h017D;    16'd27090: out <= 16'h040D;    16'd27091: out <= 16'hFD8F;
    16'd27092: out <= 16'h098F;    16'd27093: out <= 16'h0A81;    16'd27094: out <= 16'h0CC9;    16'd27095: out <= 16'h01A5;
    16'd27096: out <= 16'h04B7;    16'd27097: out <= 16'h044E;    16'd27098: out <= 16'hFFAB;    16'd27099: out <= 16'h0382;
    16'd27100: out <= 16'h00E4;    16'd27101: out <= 16'h0080;    16'd27102: out <= 16'h0647;    16'd27103: out <= 16'hFAB3;
    16'd27104: out <= 16'h0718;    16'd27105: out <= 16'hFFB3;    16'd27106: out <= 16'hF7CA;    16'd27107: out <= 16'h0033;
    16'd27108: out <= 16'h0385;    16'd27109: out <= 16'h0123;    16'd27110: out <= 16'h01CE;    16'd27111: out <= 16'hFE24;
    16'd27112: out <= 16'hFBBA;    16'd27113: out <= 16'hF2D2;    16'd27114: out <= 16'hFBE4;    16'd27115: out <= 16'hFBA9;
    16'd27116: out <= 16'hFD92;    16'd27117: out <= 16'hFE9E;    16'd27118: out <= 16'h06C1;    16'd27119: out <= 16'h0099;
    16'd27120: out <= 16'hFF7A;    16'd27121: out <= 16'hFE72;    16'd27122: out <= 16'hF6C8;    16'd27123: out <= 16'hFCC8;
    16'd27124: out <= 16'hFDE1;    16'd27125: out <= 16'hFB1D;    16'd27126: out <= 16'h01E0;    16'd27127: out <= 16'hFE84;
    16'd27128: out <= 16'h00FE;    16'd27129: out <= 16'h012A;    16'd27130: out <= 16'hFED0;    16'd27131: out <= 16'hFE52;
    16'd27132: out <= 16'hFEA3;    16'd27133: out <= 16'h0260;    16'd27134: out <= 16'hFA35;    16'd27135: out <= 16'hFCF9;
    16'd27136: out <= 16'hF964;    16'd27137: out <= 16'hFD8E;    16'd27138: out <= 16'hFB60;    16'd27139: out <= 16'hFFC5;
    16'd27140: out <= 16'hFF45;    16'd27141: out <= 16'hFED5;    16'd27142: out <= 16'hF9EB;    16'd27143: out <= 16'hFE88;
    16'd27144: out <= 16'h03BB;    16'd27145: out <= 16'hF9F6;    16'd27146: out <= 16'h05B6;    16'd27147: out <= 16'h00F0;
    16'd27148: out <= 16'h00F9;    16'd27149: out <= 16'h009D;    16'd27150: out <= 16'h01CD;    16'd27151: out <= 16'h0095;
    16'd27152: out <= 16'hFF29;    16'd27153: out <= 16'hFA33;    16'd27154: out <= 16'hFC1C;    16'd27155: out <= 16'h0140;
    16'd27156: out <= 16'hFE3E;    16'd27157: out <= 16'h0086;    16'd27158: out <= 16'hFF85;    16'd27159: out <= 16'hFEF4;
    16'd27160: out <= 16'h011F;    16'd27161: out <= 16'hFD46;    16'd27162: out <= 16'h0162;    16'd27163: out <= 16'hFC0E;
    16'd27164: out <= 16'hFD02;    16'd27165: out <= 16'hFF3F;    16'd27166: out <= 16'hFE32;    16'd27167: out <= 16'h02F5;
    16'd27168: out <= 16'hFD58;    16'd27169: out <= 16'h0481;    16'd27170: out <= 16'hFF93;    16'd27171: out <= 16'h047E;
    16'd27172: out <= 16'h0ACE;    16'd27173: out <= 16'h01DB;    16'd27174: out <= 16'h0C01;    16'd27175: out <= 16'h0BB9;
    16'd27176: out <= 16'h0831;    16'd27177: out <= 16'hFB7A;    16'd27178: out <= 16'h02B8;    16'd27179: out <= 16'h0308;
    16'd27180: out <= 16'h0871;    16'd27181: out <= 16'h075D;    16'd27182: out <= 16'h020E;    16'd27183: out <= 16'h0498;
    16'd27184: out <= 16'h0381;    16'd27185: out <= 16'h034F;    16'd27186: out <= 16'h0574;    16'd27187: out <= 16'h0395;
    16'd27188: out <= 16'h078E;    16'd27189: out <= 16'h00A7;    16'd27190: out <= 16'hFF39;    16'd27191: out <= 16'h078A;
    16'd27192: out <= 16'h0131;    16'd27193: out <= 16'h0640;    16'd27194: out <= 16'h0651;    16'd27195: out <= 16'hFD09;
    16'd27196: out <= 16'h0419;    16'd27197: out <= 16'h02F7;    16'd27198: out <= 16'h05BF;    16'd27199: out <= 16'h020D;
    16'd27200: out <= 16'h0311;    16'd27201: out <= 16'h0204;    16'd27202: out <= 16'hFAD9;    16'd27203: out <= 16'hFEE7;
    16'd27204: out <= 16'h02F6;    16'd27205: out <= 16'h024C;    16'd27206: out <= 16'h04A9;    16'd27207: out <= 16'h0961;
    16'd27208: out <= 16'h0231;    16'd27209: out <= 16'h03C7;    16'd27210: out <= 16'h05B5;    16'd27211: out <= 16'h0084;
    16'd27212: out <= 16'h02B0;    16'd27213: out <= 16'h0642;    16'd27214: out <= 16'h00BB;    16'd27215: out <= 16'h0A38;
    16'd27216: out <= 16'h06C7;    16'd27217: out <= 16'h0BD0;    16'd27218: out <= 16'h0533;    16'd27219: out <= 16'h0585;
    16'd27220: out <= 16'h04D9;    16'd27221: out <= 16'h04A4;    16'd27222: out <= 16'h04EC;    16'd27223: out <= 16'h0067;
    16'd27224: out <= 16'h0191;    16'd27225: out <= 16'h0280;    16'd27226: out <= 16'hFE8F;    16'd27227: out <= 16'h0938;
    16'd27228: out <= 16'h039A;    16'd27229: out <= 16'h02FB;    16'd27230: out <= 16'h0237;    16'd27231: out <= 16'h040F;
    16'd27232: out <= 16'h03EE;    16'd27233: out <= 16'hFEE2;    16'd27234: out <= 16'h040D;    16'd27235: out <= 16'h00F6;
    16'd27236: out <= 16'h0D01;    16'd27237: out <= 16'hFE05;    16'd27238: out <= 16'hFDC2;    16'd27239: out <= 16'h0132;
    16'd27240: out <= 16'h05CD;    16'd27241: out <= 16'h02B9;    16'd27242: out <= 16'h0407;    16'd27243: out <= 16'h08BB;
    16'd27244: out <= 16'h035C;    16'd27245: out <= 16'hFA08;    16'd27246: out <= 16'h0144;    16'd27247: out <= 16'h04A7;
    16'd27248: out <= 16'hFEA5;    16'd27249: out <= 16'h0BF4;    16'd27250: out <= 16'hFF90;    16'd27251: out <= 16'hFE72;
    16'd27252: out <= 16'h05BF;    16'd27253: out <= 16'hFF28;    16'd27254: out <= 16'h04E1;    16'd27255: out <= 16'h038A;
    16'd27256: out <= 16'h0011;    16'd27257: out <= 16'h05AD;    16'd27258: out <= 16'h0BAB;    16'd27259: out <= 16'h068C;
    16'd27260: out <= 16'h0A44;    16'd27261: out <= 16'h030C;    16'd27262: out <= 16'h0273;    16'd27263: out <= 16'h035F;
    16'd27264: out <= 16'h0B9F;    16'd27265: out <= 16'h00F7;    16'd27266: out <= 16'h0260;    16'd27267: out <= 16'h0062;
    16'd27268: out <= 16'h09B9;    16'd27269: out <= 16'h07AE;    16'd27270: out <= 16'hFC4E;    16'd27271: out <= 16'h08EE;
    16'd27272: out <= 16'h075C;    16'd27273: out <= 16'h01B4;    16'd27274: out <= 16'h061F;    16'd27275: out <= 16'h065F;
    16'd27276: out <= 16'h0001;    16'd27277: out <= 16'h0420;    16'd27278: out <= 16'h03DB;    16'd27279: out <= 16'h0470;
    16'd27280: out <= 16'h0A1B;    16'd27281: out <= 16'h0609;    16'd27282: out <= 16'h0564;    16'd27283: out <= 16'h0478;
    16'd27284: out <= 16'h02A8;    16'd27285: out <= 16'h0513;    16'd27286: out <= 16'h05B9;    16'd27287: out <= 16'h041F;
    16'd27288: out <= 16'h0236;    16'd27289: out <= 16'h0273;    16'd27290: out <= 16'h05D6;    16'd27291: out <= 16'h03A0;
    16'd27292: out <= 16'h054B;    16'd27293: out <= 16'h0075;    16'd27294: out <= 16'h066D;    16'd27295: out <= 16'h0215;
    16'd27296: out <= 16'h09B9;    16'd27297: out <= 16'h0D6E;    16'd27298: out <= 16'h01D7;    16'd27299: out <= 16'hFAC4;
    16'd27300: out <= 16'hFB34;    16'd27301: out <= 16'h02F4;    16'd27302: out <= 16'h0188;    16'd27303: out <= 16'h0159;
    16'd27304: out <= 16'hFD95;    16'd27305: out <= 16'h0139;    16'd27306: out <= 16'hFAFD;    16'd27307: out <= 16'h04E4;
    16'd27308: out <= 16'h05F2;    16'd27309: out <= 16'h00D4;    16'd27310: out <= 16'hFCF0;    16'd27311: out <= 16'hFEDB;
    16'd27312: out <= 16'h04C2;    16'd27313: out <= 16'hFE80;    16'd27314: out <= 16'h0788;    16'd27315: out <= 16'hFE8A;
    16'd27316: out <= 16'hFE8B;    16'd27317: out <= 16'h018C;    16'd27318: out <= 16'h0617;    16'd27319: out <= 16'hFFDD;
    16'd27320: out <= 16'hFE8F;    16'd27321: out <= 16'h03CA;    16'd27322: out <= 16'h07D0;    16'd27323: out <= 16'h0477;
    16'd27324: out <= 16'hFD75;    16'd27325: out <= 16'h00AE;    16'd27326: out <= 16'h054E;    16'd27327: out <= 16'h04A9;
    16'd27328: out <= 16'h0295;    16'd27329: out <= 16'hFE5B;    16'd27330: out <= 16'h0405;    16'd27331: out <= 16'h02E9;
    16'd27332: out <= 16'h024E;    16'd27333: out <= 16'hFDFA;    16'd27334: out <= 16'h0B5B;    16'd27335: out <= 16'h0476;
    16'd27336: out <= 16'hFCDA;    16'd27337: out <= 16'h0283;    16'd27338: out <= 16'h0057;    16'd27339: out <= 16'h02B0;
    16'd27340: out <= 16'h0847;    16'd27341: out <= 16'h08D3;    16'd27342: out <= 16'h0696;    16'd27343: out <= 16'h0381;
    16'd27344: out <= 16'h03FE;    16'd27345: out <= 16'hFE36;    16'd27346: out <= 16'h0564;    16'd27347: out <= 16'h025D;
    16'd27348: out <= 16'h08A9;    16'd27349: out <= 16'h03DA;    16'd27350: out <= 16'h0679;    16'd27351: out <= 16'h006F;
    16'd27352: out <= 16'hFE41;    16'd27353: out <= 16'hFC18;    16'd27354: out <= 16'h01D7;    16'd27355: out <= 16'hF342;
    16'd27356: out <= 16'hFFB4;    16'd27357: out <= 16'h0110;    16'd27358: out <= 16'hFEF7;    16'd27359: out <= 16'hFF5D;
    16'd27360: out <= 16'hFF25;    16'd27361: out <= 16'hFFA0;    16'd27362: out <= 16'hFF39;    16'd27363: out <= 16'h0074;
    16'd27364: out <= 16'hFB1C;    16'd27365: out <= 16'hFC80;    16'd27366: out <= 16'h0246;    16'd27367: out <= 16'h09BC;
    16'd27368: out <= 16'hFD75;    16'd27369: out <= 16'h05C5;    16'd27370: out <= 16'h0013;    16'd27371: out <= 16'h02FA;
    16'd27372: out <= 16'h00B2;    16'd27373: out <= 16'hFEDC;    16'd27374: out <= 16'h0090;    16'd27375: out <= 16'hFEDF;
    16'd27376: out <= 16'hFBF0;    16'd27377: out <= 16'hFDC0;    16'd27378: out <= 16'h049E;    16'd27379: out <= 16'hF6D1;
    16'd27380: out <= 16'h03AD;    16'd27381: out <= 16'hFB69;    16'd27382: out <= 16'h0342;    16'd27383: out <= 16'h01DC;
    16'd27384: out <= 16'h021A;    16'd27385: out <= 16'hFED0;    16'd27386: out <= 16'h086F;    16'd27387: out <= 16'hFDF7;
    16'd27388: out <= 16'h0106;    16'd27389: out <= 16'h02F6;    16'd27390: out <= 16'h02D5;    16'd27391: out <= 16'h0294;
    16'd27392: out <= 16'h0491;    16'd27393: out <= 16'hFACC;    16'd27394: out <= 16'h041C;    16'd27395: out <= 16'h021D;
    16'd27396: out <= 16'hFE01;    16'd27397: out <= 16'h02E1;    16'd27398: out <= 16'h064C;    16'd27399: out <= 16'h059E;
    16'd27400: out <= 16'hFF58;    16'd27401: out <= 16'h06FD;    16'd27402: out <= 16'h03C9;    16'd27403: out <= 16'hFE76;
    16'd27404: out <= 16'h0353;    16'd27405: out <= 16'h0331;    16'd27406: out <= 16'h01A1;    16'd27407: out <= 16'h0402;
    16'd27408: out <= 16'hFF56;    16'd27409: out <= 16'h02A6;    16'd27410: out <= 16'hFB9B;    16'd27411: out <= 16'hF7D3;
    16'd27412: out <= 16'hFFA0;    16'd27413: out <= 16'h08BC;    16'd27414: out <= 16'h025D;    16'd27415: out <= 16'h03D2;
    16'd27416: out <= 16'h0114;    16'd27417: out <= 16'h0161;    16'd27418: out <= 16'h0190;    16'd27419: out <= 16'h02F8;
    16'd27420: out <= 16'hFDF1;    16'd27421: out <= 16'hFF14;    16'd27422: out <= 16'hFE1A;    16'd27423: out <= 16'h0459;
    16'd27424: out <= 16'hFEE0;    16'd27425: out <= 16'h072B;    16'd27426: out <= 16'h0B56;    16'd27427: out <= 16'h0623;
    16'd27428: out <= 16'h0270;    16'd27429: out <= 16'h0C42;    16'd27430: out <= 16'h0888;    16'd27431: out <= 16'h00DF;
    16'd27432: out <= 16'h001F;    16'd27433: out <= 16'h075A;    16'd27434: out <= 16'h02AE;    16'd27435: out <= 16'h078D;
    16'd27436: out <= 16'h05B6;    16'd27437: out <= 16'h02BA;    16'd27438: out <= 16'hFFA5;    16'd27439: out <= 16'h038B;
    16'd27440: out <= 16'h01AB;    16'd27441: out <= 16'h0569;    16'd27442: out <= 16'h06E9;    16'd27443: out <= 16'h03F1;
    16'd27444: out <= 16'h0AA5;    16'd27445: out <= 16'h024F;    16'd27446: out <= 16'h09CF;    16'd27447: out <= 16'hFBD8;
    16'd27448: out <= 16'h04C9;    16'd27449: out <= 16'h01F4;    16'd27450: out <= 16'h004F;    16'd27451: out <= 16'h07EB;
    16'd27452: out <= 16'h015D;    16'd27453: out <= 16'h0CC8;    16'd27454: out <= 16'h0643;    16'd27455: out <= 16'h05B0;
    16'd27456: out <= 16'h0368;    16'd27457: out <= 16'h0465;    16'd27458: out <= 16'h032D;    16'd27459: out <= 16'h0486;
    16'd27460: out <= 16'hFFAA;    16'd27461: out <= 16'h0325;    16'd27462: out <= 16'h0521;    16'd27463: out <= 16'h0995;
    16'd27464: out <= 16'hFF7C;    16'd27465: out <= 16'h06C5;    16'd27466: out <= 16'h05CA;    16'd27467: out <= 16'h0185;
    16'd27468: out <= 16'hFCB7;    16'd27469: out <= 16'h031D;    16'd27470: out <= 16'h0112;    16'd27471: out <= 16'h0A7E;
    16'd27472: out <= 16'h038E;    16'd27473: out <= 16'h03C1;    16'd27474: out <= 16'hFE35;    16'd27475: out <= 16'h0422;
    16'd27476: out <= 16'h05A5;    16'd27477: out <= 16'h0349;    16'd27478: out <= 16'h0758;    16'd27479: out <= 16'h06DC;
    16'd27480: out <= 16'h0725;    16'd27481: out <= 16'h01F2;    16'd27482: out <= 16'h0B7F;    16'd27483: out <= 16'h0725;
    16'd27484: out <= 16'h0364;    16'd27485: out <= 16'h04E9;    16'd27486: out <= 16'h02D7;    16'd27487: out <= 16'h0577;
    16'd27488: out <= 16'h0271;    16'd27489: out <= 16'h066E;    16'd27490: out <= 16'h03D4;    16'd27491: out <= 16'hFEC6;
    16'd27492: out <= 16'h07CB;    16'd27493: out <= 16'h04E6;    16'd27494: out <= 16'h077E;    16'd27495: out <= 16'h040A;
    16'd27496: out <= 16'h0515;    16'd27497: out <= 16'h057B;    16'd27498: out <= 16'h04C4;    16'd27499: out <= 16'h0144;
    16'd27500: out <= 16'h02B4;    16'd27501: out <= 16'h03CF;    16'd27502: out <= 16'h04E5;    16'd27503: out <= 16'h01A5;
    16'd27504: out <= 16'h0C4F;    16'd27505: out <= 16'h003D;    16'd27506: out <= 16'h0956;    16'd27507: out <= 16'h03BA;
    16'd27508: out <= 16'hFF3C;    16'd27509: out <= 16'h0806;    16'd27510: out <= 16'h036C;    16'd27511: out <= 16'h0330;
    16'd27512: out <= 16'h0A84;    16'd27513: out <= 16'hFF18;    16'd27514: out <= 16'h0B59;    16'd27515: out <= 16'h072A;
    16'd27516: out <= 16'h0667;    16'd27517: out <= 16'h09CD;    16'd27518: out <= 16'h0954;    16'd27519: out <= 16'hFBB1;
    16'd27520: out <= 16'h0505;    16'd27521: out <= 16'h03D8;    16'd27522: out <= 16'hFC76;    16'd27523: out <= 16'hFF39;
    16'd27524: out <= 16'h0582;    16'd27525: out <= 16'hFF65;    16'd27526: out <= 16'h0377;    16'd27527: out <= 16'h0408;
    16'd27528: out <= 16'h05C3;    16'd27529: out <= 16'h02DD;    16'd27530: out <= 16'h006B;    16'd27531: out <= 16'hFC3E;
    16'd27532: out <= 16'h0158;    16'd27533: out <= 16'h0CC4;    16'd27534: out <= 16'h05C0;    16'd27535: out <= 16'h0555;
    16'd27536: out <= 16'h094A;    16'd27537: out <= 16'h043F;    16'd27538: out <= 16'h029B;    16'd27539: out <= 16'h0473;
    16'd27540: out <= 16'h000A;    16'd27541: out <= 16'h04B7;    16'd27542: out <= 16'hFFFF;    16'd27543: out <= 16'h0824;
    16'd27544: out <= 16'h0535;    16'd27545: out <= 16'h0008;    16'd27546: out <= 16'h0766;    16'd27547: out <= 16'h0402;
    16'd27548: out <= 16'h0078;    16'd27549: out <= 16'h03F6;    16'd27550: out <= 16'h0550;    16'd27551: out <= 16'h0415;
    16'd27552: out <= 16'h06AF;    16'd27553: out <= 16'h02C1;    16'd27554: out <= 16'h04FA;    16'd27555: out <= 16'h03B0;
    16'd27556: out <= 16'h05C1;    16'd27557: out <= 16'h0411;    16'd27558: out <= 16'hFB91;    16'd27559: out <= 16'h000D;
    16'd27560: out <= 16'hFF16;    16'd27561: out <= 16'h02C4;    16'd27562: out <= 16'h04D0;    16'd27563: out <= 16'h0319;
    16'd27564: out <= 16'h0171;    16'd27565: out <= 16'h0878;    16'd27566: out <= 16'h00DC;    16'd27567: out <= 16'h0109;
    16'd27568: out <= 16'h029C;    16'd27569: out <= 16'h0389;    16'd27570: out <= 16'h032F;    16'd27571: out <= 16'h0229;
    16'd27572: out <= 16'hFBE9;    16'd27573: out <= 16'h0086;    16'd27574: out <= 16'hFC28;    16'd27575: out <= 16'h02F8;
    16'd27576: out <= 16'hF8D3;    16'd27577: out <= 16'h0EA2;    16'd27578: out <= 16'h065B;    16'd27579: out <= 16'h047A;
    16'd27580: out <= 16'h06C0;    16'd27581: out <= 16'h03F9;    16'd27582: out <= 16'hFE07;    16'd27583: out <= 16'h0159;
    16'd27584: out <= 16'h0036;    16'd27585: out <= 16'hFEBD;    16'd27586: out <= 16'hFFCF;    16'd27587: out <= 16'h0918;
    16'd27588: out <= 16'h0571;    16'd27589: out <= 16'h0241;    16'd27590: out <= 16'h0369;    16'd27591: out <= 16'h08F0;
    16'd27592: out <= 16'h0361;    16'd27593: out <= 16'h08CE;    16'd27594: out <= 16'h029E;    16'd27595: out <= 16'h06D3;
    16'd27596: out <= 16'hFEC2;    16'd27597: out <= 16'h0570;    16'd27598: out <= 16'h033B;    16'd27599: out <= 16'h06D3;
    16'd27600: out <= 16'h0273;    16'd27601: out <= 16'hFEFB;    16'd27602: out <= 16'hFDC3;    16'd27603: out <= 16'h017A;
    16'd27604: out <= 16'hFF87;    16'd27605: out <= 16'h0447;    16'd27606: out <= 16'h03F7;    16'd27607: out <= 16'h0009;
    16'd27608: out <= 16'h08A6;    16'd27609: out <= 16'h0500;    16'd27610: out <= 16'hFF78;    16'd27611: out <= 16'hFB58;
    16'd27612: out <= 16'h02EA;    16'd27613: out <= 16'h0252;    16'd27614: out <= 16'hFF0C;    16'd27615: out <= 16'h0040;
    16'd27616: out <= 16'hFD9C;    16'd27617: out <= 16'hFC63;    16'd27618: out <= 16'h02AE;    16'd27619: out <= 16'hF9F1;
    16'd27620: out <= 16'h056C;    16'd27621: out <= 16'h00C5;    16'd27622: out <= 16'h0012;    16'd27623: out <= 16'hFD4F;
    16'd27624: out <= 16'h0180;    16'd27625: out <= 16'h0299;    16'd27626: out <= 16'hFA80;    16'd27627: out <= 16'h0108;
    16'd27628: out <= 16'h024B;    16'd27629: out <= 16'hFECF;    16'd27630: out <= 16'h0246;    16'd27631: out <= 16'h0276;
    16'd27632: out <= 16'hFF98;    16'd27633: out <= 16'h0118;    16'd27634: out <= 16'h09C3;    16'd27635: out <= 16'hFDE8;
    16'd27636: out <= 16'h0110;    16'd27637: out <= 16'h02C4;    16'd27638: out <= 16'h02A5;    16'd27639: out <= 16'h02B3;
    16'd27640: out <= 16'hFB79;    16'd27641: out <= 16'h00FC;    16'd27642: out <= 16'hFB20;    16'd27643: out <= 16'h0612;
    16'd27644: out <= 16'h0749;    16'd27645: out <= 16'h01D2;    16'd27646: out <= 16'h0652;    16'd27647: out <= 16'h004D;
    16'd27648: out <= 16'h066D;    16'd27649: out <= 16'h063B;    16'd27650: out <= 16'hFDA3;    16'd27651: out <= 16'h0328;
    16'd27652: out <= 16'hFD51;    16'd27653: out <= 16'h035D;    16'd27654: out <= 16'h006F;    16'd27655: out <= 16'hFD1D;
    16'd27656: out <= 16'hFB4B;    16'd27657: out <= 16'h006A;    16'd27658: out <= 16'hFC29;    16'd27659: out <= 16'h0944;
    16'd27660: out <= 16'h01FD;    16'd27661: out <= 16'h00F0;    16'd27662: out <= 16'h0050;    16'd27663: out <= 16'hFAFF;
    16'd27664: out <= 16'hFE3D;    16'd27665: out <= 16'h01BF;    16'd27666: out <= 16'h032F;    16'd27667: out <= 16'h044F;
    16'd27668: out <= 16'h04C0;    16'd27669: out <= 16'h0423;    16'd27670: out <= 16'h0871;    16'd27671: out <= 16'hFBB3;
    16'd27672: out <= 16'h07F4;    16'd27673: out <= 16'h0527;    16'd27674: out <= 16'hF399;    16'd27675: out <= 16'h043B;
    16'd27676: out <= 16'hFFC4;    16'd27677: out <= 16'h0CF7;    16'd27678: out <= 16'h020B;    16'd27679: out <= 16'hF938;
    16'd27680: out <= 16'hFEF4;    16'd27681: out <= 16'h00E8;    16'd27682: out <= 16'h0391;    16'd27683: out <= 16'h0264;
    16'd27684: out <= 16'h0CEB;    16'd27685: out <= 16'h0191;    16'd27686: out <= 16'h033D;    16'd27687: out <= 16'h0476;
    16'd27688: out <= 16'h04B1;    16'd27689: out <= 16'h0682;    16'd27690: out <= 16'hFE5A;    16'd27691: out <= 16'h091B;
    16'd27692: out <= 16'h0346;    16'd27693: out <= 16'h0A91;    16'd27694: out <= 16'h07D6;    16'd27695: out <= 16'h061E;
    16'd27696: out <= 16'h03BE;    16'd27697: out <= 16'h00DE;    16'd27698: out <= 16'hFFF7;    16'd27699: out <= 16'h01BA;
    16'd27700: out <= 16'h001A;    16'd27701: out <= 16'hFF71;    16'd27702: out <= 16'h0699;    16'd27703: out <= 16'h083B;
    16'd27704: out <= 16'h0604;    16'd27705: out <= 16'h093E;    16'd27706: out <= 16'h0220;    16'd27707: out <= 16'h0B93;
    16'd27708: out <= 16'h064E;    16'd27709: out <= 16'h0C10;    16'd27710: out <= 16'h04DB;    16'd27711: out <= 16'h061A;
    16'd27712: out <= 16'h069A;    16'd27713: out <= 16'h03FC;    16'd27714: out <= 16'h0832;    16'd27715: out <= 16'hFF4E;
    16'd27716: out <= 16'h08B0;    16'd27717: out <= 16'hFD83;    16'd27718: out <= 16'h0606;    16'd27719: out <= 16'h06A0;
    16'd27720: out <= 16'hFF85;    16'd27721: out <= 16'h0193;    16'd27722: out <= 16'h076A;    16'd27723: out <= 16'h0060;
    16'd27724: out <= 16'hFFDF;    16'd27725: out <= 16'h04AA;    16'd27726: out <= 16'h0524;    16'd27727: out <= 16'h0B81;
    16'd27728: out <= 16'h04C6;    16'd27729: out <= 16'h068C;    16'd27730: out <= 16'h0089;    16'd27731: out <= 16'h0161;
    16'd27732: out <= 16'h0981;    16'd27733: out <= 16'h0131;    16'd27734: out <= 16'hFF1D;    16'd27735: out <= 16'h0562;
    16'd27736: out <= 16'h0404;    16'd27737: out <= 16'h0BBF;    16'd27738: out <= 16'h039E;    16'd27739: out <= 16'h06D2;
    16'd27740: out <= 16'hFCFE;    16'd27741: out <= 16'h0010;    16'd27742: out <= 16'hFCF7;    16'd27743: out <= 16'h07A2;
    16'd27744: out <= 16'h0960;    16'd27745: out <= 16'h0238;    16'd27746: out <= 16'h04DD;    16'd27747: out <= 16'h03E0;
    16'd27748: out <= 16'h02AC;    16'd27749: out <= 16'h0249;    16'd27750: out <= 16'h0A64;    16'd27751: out <= 16'h090C;
    16'd27752: out <= 16'h0770;    16'd27753: out <= 16'hFFF5;    16'd27754: out <= 16'h063B;    16'd27755: out <= 16'h041F;
    16'd27756: out <= 16'h0510;    16'd27757: out <= 16'h023D;    16'd27758: out <= 16'h0340;    16'd27759: out <= 16'h03B3;
    16'd27760: out <= 16'h049B;    16'd27761: out <= 16'h0261;    16'd27762: out <= 16'hFDF6;    16'd27763: out <= 16'h04EF;
    16'd27764: out <= 16'h0721;    16'd27765: out <= 16'h0717;    16'd27766: out <= 16'h060D;    16'd27767: out <= 16'h09F0;
    16'd27768: out <= 16'h0494;    16'd27769: out <= 16'h03A8;    16'd27770: out <= 16'h065E;    16'd27771: out <= 16'h05CF;
    16'd27772: out <= 16'h0850;    16'd27773: out <= 16'h05D6;    16'd27774: out <= 16'h0810;    16'd27775: out <= 16'h01BD;
    16'd27776: out <= 16'h0298;    16'd27777: out <= 16'hFE07;    16'd27778: out <= 16'hFF17;    16'd27779: out <= 16'h04A1;
    16'd27780: out <= 16'h02AA;    16'd27781: out <= 16'h008A;    16'd27782: out <= 16'h04F2;    16'd27783: out <= 16'h009A;
    16'd27784: out <= 16'h01EB;    16'd27785: out <= 16'h0874;    16'd27786: out <= 16'h0694;    16'd27787: out <= 16'h02C3;
    16'd27788: out <= 16'h04F0;    16'd27789: out <= 16'h05A9;    16'd27790: out <= 16'h0403;    16'd27791: out <= 16'h08F3;
    16'd27792: out <= 16'h01E2;    16'd27793: out <= 16'hFFB0;    16'd27794: out <= 16'h0385;    16'd27795: out <= 16'h07EA;
    16'd27796: out <= 16'h022A;    16'd27797: out <= 16'h02DA;    16'd27798: out <= 16'h0289;    16'd27799: out <= 16'h02E4;
    16'd27800: out <= 16'h0851;    16'd27801: out <= 16'h05B1;    16'd27802: out <= 16'h01F3;    16'd27803: out <= 16'h0383;
    16'd27804: out <= 16'h03D5;    16'd27805: out <= 16'h0639;    16'd27806: out <= 16'h00B7;    16'd27807: out <= 16'h0460;
    16'd27808: out <= 16'h0461;    16'd27809: out <= 16'h08C8;    16'd27810: out <= 16'h0591;    16'd27811: out <= 16'h06D6;
    16'd27812: out <= 16'hFFA2;    16'd27813: out <= 16'hFD4F;    16'd27814: out <= 16'h09E6;    16'd27815: out <= 16'hFE05;
    16'd27816: out <= 16'h070E;    16'd27817: out <= 16'h0352;    16'd27818: out <= 16'h0A3E;    16'd27819: out <= 16'h0791;
    16'd27820: out <= 16'h0306;    16'd27821: out <= 16'h0114;    16'd27822: out <= 16'h063E;    16'd27823: out <= 16'h094A;
    16'd27824: out <= 16'h08F7;    16'd27825: out <= 16'h0803;    16'd27826: out <= 16'h0244;    16'd27827: out <= 16'h05A0;
    16'd27828: out <= 16'h09B5;    16'd27829: out <= 16'hF8ED;    16'd27830: out <= 16'hFC2A;    16'd27831: out <= 16'hFFC1;
    16'd27832: out <= 16'hFF1C;    16'd27833: out <= 16'h00A1;    16'd27834: out <= 16'h04FE;    16'd27835: out <= 16'h0028;
    16'd27836: out <= 16'hFED8;    16'd27837: out <= 16'h091A;    16'd27838: out <= 16'hFE9B;    16'd27839: out <= 16'hFB64;
    16'd27840: out <= 16'h080B;    16'd27841: out <= 16'h03B8;    16'd27842: out <= 16'h07E6;    16'd27843: out <= 16'h0A86;
    16'd27844: out <= 16'h04C4;    16'd27845: out <= 16'h02C9;    16'd27846: out <= 16'hFF63;    16'd27847: out <= 16'h0427;
    16'd27848: out <= 16'h0272;    16'd27849: out <= 16'h0868;    16'd27850: out <= 16'h0425;    16'd27851: out <= 16'h0A64;
    16'd27852: out <= 16'h0607;    16'd27853: out <= 16'hFE80;    16'd27854: out <= 16'h05D7;    16'd27855: out <= 16'h0225;
    16'd27856: out <= 16'h01E6;    16'd27857: out <= 16'h087C;    16'd27858: out <= 16'h0731;    16'd27859: out <= 16'h033A;
    16'd27860: out <= 16'hFF05;    16'd27861: out <= 16'h0220;    16'd27862: out <= 16'hFEA1;    16'd27863: out <= 16'h0186;
    16'd27864: out <= 16'h0115;    16'd27865: out <= 16'h02E6;    16'd27866: out <= 16'h04F5;    16'd27867: out <= 16'hFC22;
    16'd27868: out <= 16'h00CF;    16'd27869: out <= 16'h02D0;    16'd27870: out <= 16'h04D7;    16'd27871: out <= 16'h0027;
    16'd27872: out <= 16'hFCAD;    16'd27873: out <= 16'h0A6A;    16'd27874: out <= 16'h05E3;    16'd27875: out <= 16'hFE3D;
    16'd27876: out <= 16'h01DD;    16'd27877: out <= 16'h03EF;    16'd27878: out <= 16'h040B;    16'd27879: out <= 16'hFA88;
    16'd27880: out <= 16'hFE8E;    16'd27881: out <= 16'hFC7B;    16'd27882: out <= 16'hFC1D;    16'd27883: out <= 16'h00E6;
    16'd27884: out <= 16'hF9D8;    16'd27885: out <= 16'h074A;    16'd27886: out <= 16'hFDA0;    16'd27887: out <= 16'h0862;
    16'd27888: out <= 16'hFE35;    16'd27889: out <= 16'h01F8;    16'd27890: out <= 16'h0089;    16'd27891: out <= 16'h0578;
    16'd27892: out <= 16'hFFAE;    16'd27893: out <= 16'hFA76;    16'd27894: out <= 16'h03D8;    16'd27895: out <= 16'hFA1A;
    16'd27896: out <= 16'h00F7;    16'd27897: out <= 16'hFFA1;    16'd27898: out <= 16'h0002;    16'd27899: out <= 16'h0198;
    16'd27900: out <= 16'h01F3;    16'd27901: out <= 16'h07FC;    16'd27902: out <= 16'hF96F;    16'd27903: out <= 16'hFF53;
    16'd27904: out <= 16'h0421;    16'd27905: out <= 16'hFFF2;    16'd27906: out <= 16'h0360;    16'd27907: out <= 16'h097B;
    16'd27908: out <= 16'hFDC8;    16'd27909: out <= 16'h0606;    16'd27910: out <= 16'h0603;    16'd27911: out <= 16'hFAB3;
    16'd27912: out <= 16'h0818;    16'd27913: out <= 16'hFDB5;    16'd27914: out <= 16'h0470;    16'd27915: out <= 16'hFD33;
    16'd27916: out <= 16'hFFAB;    16'd27917: out <= 16'h017E;    16'd27918: out <= 16'h00FB;    16'd27919: out <= 16'h0296;
    16'd27920: out <= 16'hFAFA;    16'd27921: out <= 16'h03C9;    16'd27922: out <= 16'h03FB;    16'd27923: out <= 16'h004F;
    16'd27924: out <= 16'hFECB;    16'd27925: out <= 16'h043F;    16'd27926: out <= 16'hFC8E;    16'd27927: out <= 16'h0136;
    16'd27928: out <= 16'h036A;    16'd27929: out <= 16'h00A7;    16'd27930: out <= 16'h0471;    16'd27931: out <= 16'h03D8;
    16'd27932: out <= 16'h0609;    16'd27933: out <= 16'hFCBE;    16'd27934: out <= 16'h03C7;    16'd27935: out <= 16'h0120;
    16'd27936: out <= 16'h026A;    16'd27937: out <= 16'h0332;    16'd27938: out <= 16'h019A;    16'd27939: out <= 16'h0730;
    16'd27940: out <= 16'h0509;    16'd27941: out <= 16'h0370;    16'd27942: out <= 16'h06AA;    16'd27943: out <= 16'h04D9;
    16'd27944: out <= 16'h06DB;    16'd27945: out <= 16'hFFDF;    16'd27946: out <= 16'h0757;    16'd27947: out <= 16'h041B;
    16'd27948: out <= 16'h007D;    16'd27949: out <= 16'h03D6;    16'd27950: out <= 16'hF865;    16'd27951: out <= 16'h0322;
    16'd27952: out <= 16'h0B92;    16'd27953: out <= 16'hFDC8;    16'd27954: out <= 16'hFD42;    16'd27955: out <= 16'h0416;
    16'd27956: out <= 16'h045A;    16'd27957: out <= 16'h026A;    16'd27958: out <= 16'hFF10;    16'd27959: out <= 16'h0050;
    16'd27960: out <= 16'hFEBF;    16'd27961: out <= 16'h07C7;    16'd27962: out <= 16'h0059;    16'd27963: out <= 16'h01C7;
    16'd27964: out <= 16'h01AA;    16'd27965: out <= 16'h0582;    16'd27966: out <= 16'h033C;    16'd27967: out <= 16'hFC2D;
    16'd27968: out <= 16'h0583;    16'd27969: out <= 16'h05DC;    16'd27970: out <= 16'h057D;    16'd27971: out <= 16'h038B;
    16'd27972: out <= 16'h054E;    16'd27973: out <= 16'h037B;    16'd27974: out <= 16'h03E4;    16'd27975: out <= 16'h002B;
    16'd27976: out <= 16'h0760;    16'd27977: out <= 16'h07E7;    16'd27978: out <= 16'h02A6;    16'd27979: out <= 16'h054F;
    16'd27980: out <= 16'h0958;    16'd27981: out <= 16'h00F5;    16'd27982: out <= 16'h0647;    16'd27983: out <= 16'h0761;
    16'd27984: out <= 16'h086C;    16'd27985: out <= 16'h0BA8;    16'd27986: out <= 16'h061B;    16'd27987: out <= 16'h0426;
    16'd27988: out <= 16'h0156;    16'd27989: out <= 16'hFF2D;    16'd27990: out <= 16'h0374;    16'd27991: out <= 16'h050E;
    16'd27992: out <= 16'h00D1;    16'd27993: out <= 16'h0705;    16'd27994: out <= 16'h021D;    16'd27995: out <= 16'h088E;
    16'd27996: out <= 16'h0493;    16'd27997: out <= 16'hFFBE;    16'd27998: out <= 16'h0DC9;    16'd27999: out <= 16'h0436;
    16'd28000: out <= 16'h0172;    16'd28001: out <= 16'h02A3;    16'd28002: out <= 16'h02E7;    16'd28003: out <= 16'hF99D;
    16'd28004: out <= 16'h0581;    16'd28005: out <= 16'h0745;    16'd28006: out <= 16'hFFF0;    16'd28007: out <= 16'h09BE;
    16'd28008: out <= 16'hFC63;    16'd28009: out <= 16'h0451;    16'd28010: out <= 16'h05D2;    16'd28011: out <= 16'h01C4;
    16'd28012: out <= 16'h05E8;    16'd28013: out <= 16'h04C9;    16'd28014: out <= 16'h00F5;    16'd28015: out <= 16'hFF00;
    16'd28016: out <= 16'h0597;    16'd28017: out <= 16'h0303;    16'd28018: out <= 16'h0189;    16'd28019: out <= 16'h0038;
    16'd28020: out <= 16'h07FF;    16'd28021: out <= 16'h0994;    16'd28022: out <= 16'hFE3C;    16'd28023: out <= 16'h089B;
    16'd28024: out <= 16'h0527;    16'd28025: out <= 16'h01E5;    16'd28026: out <= 16'hFE98;    16'd28027: out <= 16'hFF39;
    16'd28028: out <= 16'h06DF;    16'd28029: out <= 16'h0A27;    16'd28030: out <= 16'h04A1;    16'd28031: out <= 16'h0D26;
    16'd28032: out <= 16'h041C;    16'd28033: out <= 16'h0671;    16'd28034: out <= 16'h05C4;    16'd28035: out <= 16'h0417;
    16'd28036: out <= 16'h0231;    16'd28037: out <= 16'hFDB3;    16'd28038: out <= 16'h06D8;    16'd28039: out <= 16'h01B9;
    16'd28040: out <= 16'h079E;    16'd28041: out <= 16'h0694;    16'd28042: out <= 16'h0B78;    16'd28043: out <= 16'h08EF;
    16'd28044: out <= 16'h0033;    16'd28045: out <= 16'h0478;    16'd28046: out <= 16'h030A;    16'd28047: out <= 16'h059F;
    16'd28048: out <= 16'h0605;    16'd28049: out <= 16'h0359;    16'd28050: out <= 16'hFFD5;    16'd28051: out <= 16'h04EA;
    16'd28052: out <= 16'h004C;    16'd28053: out <= 16'h03D3;    16'd28054: out <= 16'hFE00;    16'd28055: out <= 16'h0B16;
    16'd28056: out <= 16'h0787;    16'd28057: out <= 16'h0264;    16'd28058: out <= 16'h0513;    16'd28059: out <= 16'h0188;
    16'd28060: out <= 16'h02B0;    16'd28061: out <= 16'h0615;    16'd28062: out <= 16'h05AD;    16'd28063: out <= 16'h0731;
    16'd28064: out <= 16'h02D3;    16'd28065: out <= 16'h06C5;    16'd28066: out <= 16'h0B8D;    16'd28067: out <= 16'h03CE;
    16'd28068: out <= 16'h0431;    16'd28069: out <= 16'h0330;    16'd28070: out <= 16'hFE73;    16'd28071: out <= 16'h0961;
    16'd28072: out <= 16'hFD70;    16'd28073: out <= 16'h0607;    16'd28074: out <= 16'hF957;    16'd28075: out <= 16'hFE98;
    16'd28076: out <= 16'h0473;    16'd28077: out <= 16'h091E;    16'd28078: out <= 16'h0538;    16'd28079: out <= 16'h06F7;
    16'd28080: out <= 16'h0279;    16'd28081: out <= 16'h01C1;    16'd28082: out <= 16'h01C3;    16'd28083: out <= 16'h06FC;
    16'd28084: out <= 16'hFE51;    16'd28085: out <= 16'hFF0D;    16'd28086: out <= 16'h0031;    16'd28087: out <= 16'h0135;
    16'd28088: out <= 16'h04CB;    16'd28089: out <= 16'h009B;    16'd28090: out <= 16'h049A;    16'd28091: out <= 16'h0760;
    16'd28092: out <= 16'h0683;    16'd28093: out <= 16'h088E;    16'd28094: out <= 16'h03A0;    16'd28095: out <= 16'h03C2;
    16'd28096: out <= 16'h06EF;    16'd28097: out <= 16'h0AE8;    16'd28098: out <= 16'h063B;    16'd28099: out <= 16'h05AF;
    16'd28100: out <= 16'h0A20;    16'd28101: out <= 16'h07C7;    16'd28102: out <= 16'h0307;    16'd28103: out <= 16'h017E;
    16'd28104: out <= 16'h00C3;    16'd28105: out <= 16'h084B;    16'd28106: out <= 16'h0A5E;    16'd28107: out <= 16'h0210;
    16'd28108: out <= 16'h02C9;    16'd28109: out <= 16'h0462;    16'd28110: out <= 16'h04B4;    16'd28111: out <= 16'hFDEB;
    16'd28112: out <= 16'h08E0;    16'd28113: out <= 16'h0C4F;    16'd28114: out <= 16'h08B6;    16'd28115: out <= 16'h080B;
    16'd28116: out <= 16'h0507;    16'd28117: out <= 16'h0377;    16'd28118: out <= 16'h0256;    16'd28119: out <= 16'h06FD;
    16'd28120: out <= 16'h00EB;    16'd28121: out <= 16'h00E4;    16'd28122: out <= 16'h0134;    16'd28123: out <= 16'hF981;
    16'd28124: out <= 16'h02C8;    16'd28125: out <= 16'h046C;    16'd28126: out <= 16'h01E0;    16'd28127: out <= 16'h03F9;
    16'd28128: out <= 16'hFD3B;    16'd28129: out <= 16'h02FB;    16'd28130: out <= 16'h0A97;    16'd28131: out <= 16'h03E5;
    16'd28132: out <= 16'h04CA;    16'd28133: out <= 16'hFC0D;    16'd28134: out <= 16'hFFBF;    16'd28135: out <= 16'hFA20;
    16'd28136: out <= 16'hFC57;    16'd28137: out <= 16'h0001;    16'd28138: out <= 16'h0351;    16'd28139: out <= 16'hFCBA;
    16'd28140: out <= 16'hFF0D;    16'd28141: out <= 16'hFE3C;    16'd28142: out <= 16'hFC92;    16'd28143: out <= 16'h058E;
    16'd28144: out <= 16'h0858;    16'd28145: out <= 16'h010D;    16'd28146: out <= 16'h049D;    16'd28147: out <= 16'hFE1D;
    16'd28148: out <= 16'h02BB;    16'd28149: out <= 16'hFB9B;    16'd28150: out <= 16'h038A;    16'd28151: out <= 16'h02C9;
    16'd28152: out <= 16'hFD3E;    16'd28153: out <= 16'h065E;    16'd28154: out <= 16'hFE24;    16'd28155: out <= 16'h05C6;
    16'd28156: out <= 16'hFD87;    16'd28157: out <= 16'h0376;    16'd28158: out <= 16'h0136;    16'd28159: out <= 16'hFC10;
    16'd28160: out <= 16'hFE19;    16'd28161: out <= 16'h03B0;    16'd28162: out <= 16'h0ACE;    16'd28163: out <= 16'h0587;
    16'd28164: out <= 16'hF9CD;    16'd28165: out <= 16'h0313;    16'd28166: out <= 16'hFE7A;    16'd28167: out <= 16'h0442;
    16'd28168: out <= 16'h038E;    16'd28169: out <= 16'h013F;    16'd28170: out <= 16'hFBEB;    16'd28171: out <= 16'h05CE;
    16'd28172: out <= 16'hFF70;    16'd28173: out <= 16'h02D1;    16'd28174: out <= 16'h009B;    16'd28175: out <= 16'hFC54;
    16'd28176: out <= 16'h0484;    16'd28177: out <= 16'h0755;    16'd28178: out <= 16'h015F;    16'd28179: out <= 16'hFC9C;
    16'd28180: out <= 16'hFDE4;    16'd28181: out <= 16'h023C;    16'd28182: out <= 16'hFEB5;    16'd28183: out <= 16'h092A;
    16'd28184: out <= 16'h0587;    16'd28185: out <= 16'h0000;    16'd28186: out <= 16'h028B;    16'd28187: out <= 16'h03C4;
    16'd28188: out <= 16'h036E;    16'd28189: out <= 16'h03EF;    16'd28190: out <= 16'h0070;    16'd28191: out <= 16'h041C;
    16'd28192: out <= 16'hFB43;    16'd28193: out <= 16'h0385;    16'd28194: out <= 16'h0B74;    16'd28195: out <= 16'h06BD;
    16'd28196: out <= 16'h0AAD;    16'd28197: out <= 16'h02D8;    16'd28198: out <= 16'h030C;    16'd28199: out <= 16'hFF31;
    16'd28200: out <= 16'h0043;    16'd28201: out <= 16'h0651;    16'd28202: out <= 16'h0181;    16'd28203: out <= 16'h0648;
    16'd28204: out <= 16'h07B7;    16'd28205: out <= 16'h05CE;    16'd28206: out <= 16'h059F;    16'd28207: out <= 16'h0368;
    16'd28208: out <= 16'hFC5D;    16'd28209: out <= 16'h0B9C;    16'd28210: out <= 16'h022C;    16'd28211: out <= 16'h05EB;
    16'd28212: out <= 16'hFAD2;    16'd28213: out <= 16'h01F1;    16'd28214: out <= 16'h0608;    16'd28215: out <= 16'h005E;
    16'd28216: out <= 16'h00D0;    16'd28217: out <= 16'hFB9C;    16'd28218: out <= 16'h0077;    16'd28219: out <= 16'h04E3;
    16'd28220: out <= 16'h08D0;    16'd28221: out <= 16'h04E5;    16'd28222: out <= 16'hF9B9;    16'd28223: out <= 16'h0DF9;
    16'd28224: out <= 16'h06DD;    16'd28225: out <= 16'h055B;    16'd28226: out <= 16'h01F8;    16'd28227: out <= 16'hFD7D;
    16'd28228: out <= 16'h0A1C;    16'd28229: out <= 16'h03DF;    16'd28230: out <= 16'h0452;    16'd28231: out <= 16'h0A50;
    16'd28232: out <= 16'h0279;    16'd28233: out <= 16'h03E9;    16'd28234: out <= 16'h0351;    16'd28235: out <= 16'hFFA5;
    16'd28236: out <= 16'h0175;    16'd28237: out <= 16'h06C0;    16'd28238: out <= 16'h0360;    16'd28239: out <= 16'h04A7;
    16'd28240: out <= 16'h01F6;    16'd28241: out <= 16'h093A;    16'd28242: out <= 16'h045D;    16'd28243: out <= 16'h0447;
    16'd28244: out <= 16'h0415;    16'd28245: out <= 16'h04BC;    16'd28246: out <= 16'h02BF;    16'd28247: out <= 16'h03B6;
    16'd28248: out <= 16'h079C;    16'd28249: out <= 16'h0286;    16'd28250: out <= 16'h064D;    16'd28251: out <= 16'h02F4;
    16'd28252: out <= 16'hFD60;    16'd28253: out <= 16'h06EF;    16'd28254: out <= 16'hFF88;    16'd28255: out <= 16'h02AD;
    16'd28256: out <= 16'h083A;    16'd28257: out <= 16'h0504;    16'd28258: out <= 16'h07DE;    16'd28259: out <= 16'hFABD;
    16'd28260: out <= 16'hFF7B;    16'd28261: out <= 16'h05B5;    16'd28262: out <= 16'hFCD6;    16'd28263: out <= 16'hFD13;
    16'd28264: out <= 16'h07B0;    16'd28265: out <= 16'hFF61;    16'd28266: out <= 16'h04DD;    16'd28267: out <= 16'h078F;
    16'd28268: out <= 16'h00C2;    16'd28269: out <= 16'hFEF0;    16'd28270: out <= 16'hFFB5;    16'd28271: out <= 16'h05AD;
    16'd28272: out <= 16'hFFFB;    16'd28273: out <= 16'h0AC9;    16'd28274: out <= 16'h0411;    16'd28275: out <= 16'hFB7A;
    16'd28276: out <= 16'h0A35;    16'd28277: out <= 16'h0677;    16'd28278: out <= 16'h1061;    16'd28279: out <= 16'h093B;
    16'd28280: out <= 16'h02EA;    16'd28281: out <= 16'h049A;    16'd28282: out <= 16'h04A0;    16'd28283: out <= 16'h0519;
    16'd28284: out <= 16'h083E;    16'd28285: out <= 16'hFFF9;    16'd28286: out <= 16'hFA55;    16'd28287: out <= 16'h048E;
    16'd28288: out <= 16'h06D8;    16'd28289: out <= 16'h04D9;    16'd28290: out <= 16'h088E;    16'd28291: out <= 16'h0AD8;
    16'd28292: out <= 16'h0134;    16'd28293: out <= 16'h05D6;    16'd28294: out <= 16'h0919;    16'd28295: out <= 16'h0413;
    16'd28296: out <= 16'h049D;    16'd28297: out <= 16'h076C;    16'd28298: out <= 16'h08EF;    16'd28299: out <= 16'h0567;
    16'd28300: out <= 16'h0292;    16'd28301: out <= 16'h034E;    16'd28302: out <= 16'h0653;    16'd28303: out <= 16'h00D9;
    16'd28304: out <= 16'h0489;    16'd28305: out <= 16'h042A;    16'd28306: out <= 16'h0515;    16'd28307: out <= 16'h035D;
    16'd28308: out <= 16'h00FD;    16'd28309: out <= 16'h0969;    16'd28310: out <= 16'h0582;    16'd28311: out <= 16'h06FE;
    16'd28312: out <= 16'h05D6;    16'd28313: out <= 16'h02AF;    16'd28314: out <= 16'h039D;    16'd28315: out <= 16'h05BC;
    16'd28316: out <= 16'h03E7;    16'd28317: out <= 16'h0ADE;    16'd28318: out <= 16'h0814;    16'd28319: out <= 16'h0193;
    16'd28320: out <= 16'h08F1;    16'd28321: out <= 16'h0900;    16'd28322: out <= 16'h09CF;    16'd28323: out <= 16'h05AB;
    16'd28324: out <= 16'h0BF5;    16'd28325: out <= 16'h06A8;    16'd28326: out <= 16'h02C0;    16'd28327: out <= 16'h034D;
    16'd28328: out <= 16'h0398;    16'd28329: out <= 16'h07CD;    16'd28330: out <= 16'h02D1;    16'd28331: out <= 16'hFECB;
    16'd28332: out <= 16'h0251;    16'd28333: out <= 16'hFF1B;    16'd28334: out <= 16'hFD96;    16'd28335: out <= 16'h0249;
    16'd28336: out <= 16'h0834;    16'd28337: out <= 16'h0262;    16'd28338: out <= 16'h0493;    16'd28339: out <= 16'h0C15;
    16'd28340: out <= 16'h0222;    16'd28341: out <= 16'h005B;    16'd28342: out <= 16'h0148;    16'd28343: out <= 16'h059B;
    16'd28344: out <= 16'h0AC5;    16'd28345: out <= 16'h04F0;    16'd28346: out <= 16'h0817;    16'd28347: out <= 16'hFD01;
    16'd28348: out <= 16'h05A4;    16'd28349: out <= 16'h0074;    16'd28350: out <= 16'hFE20;    16'd28351: out <= 16'hFFDC;
    16'd28352: out <= 16'h013A;    16'd28353: out <= 16'h043F;    16'd28354: out <= 16'h0465;    16'd28355: out <= 16'h026A;
    16'd28356: out <= 16'h0992;    16'd28357: out <= 16'h0325;    16'd28358: out <= 16'h05A5;    16'd28359: out <= 16'h03A2;
    16'd28360: out <= 16'h0620;    16'd28361: out <= 16'h0B0B;    16'd28362: out <= 16'h02B8;    16'd28363: out <= 16'h074C;
    16'd28364: out <= 16'h040B;    16'd28365: out <= 16'h018D;    16'd28366: out <= 16'h0696;    16'd28367: out <= 16'h02A5;
    16'd28368: out <= 16'h0932;    16'd28369: out <= 16'h0449;    16'd28370: out <= 16'h0171;    16'd28371: out <= 16'h007A;
    16'd28372: out <= 16'h0650;    16'd28373: out <= 16'h09CF;    16'd28374: out <= 16'hFF39;    16'd28375: out <= 16'h01BB;
    16'd28376: out <= 16'h0221;    16'd28377: out <= 16'h004F;    16'd28378: out <= 16'hFE5A;    16'd28379: out <= 16'hFE06;
    16'd28380: out <= 16'h019E;    16'd28381: out <= 16'hFECA;    16'd28382: out <= 16'hFE41;    16'd28383: out <= 16'hFEFA;
    16'd28384: out <= 16'hFAC6;    16'd28385: out <= 16'hF92C;    16'd28386: out <= 16'h011E;    16'd28387: out <= 16'hFF5C;
    16'd28388: out <= 16'h00F3;    16'd28389: out <= 16'hFDAE;    16'd28390: out <= 16'hFA4D;    16'd28391: out <= 16'h01C9;
    16'd28392: out <= 16'h0130;    16'd28393: out <= 16'hFDF9;    16'd28394: out <= 16'h05FB;    16'd28395: out <= 16'h0335;
    16'd28396: out <= 16'h0045;    16'd28397: out <= 16'h018A;    16'd28398: out <= 16'h0603;    16'd28399: out <= 16'hFD16;
    16'd28400: out <= 16'hFFCE;    16'd28401: out <= 16'hFE06;    16'd28402: out <= 16'hFFC9;    16'd28403: out <= 16'h0125;
    16'd28404: out <= 16'hFF86;    16'd28405: out <= 16'hFD21;    16'd28406: out <= 16'hF5D0;    16'd28407: out <= 16'h021A;
    16'd28408: out <= 16'hFCC3;    16'd28409: out <= 16'hFDAB;    16'd28410: out <= 16'h01D6;    16'd28411: out <= 16'hFB49;
    16'd28412: out <= 16'h00FC;    16'd28413: out <= 16'hF868;    16'd28414: out <= 16'h031A;    16'd28415: out <= 16'hFAB3;
    16'd28416: out <= 16'h01FE;    16'd28417: out <= 16'h04E4;    16'd28418: out <= 16'h0369;    16'd28419: out <= 16'h03FF;
    16'd28420: out <= 16'hFEA0;    16'd28421: out <= 16'hFE68;    16'd28422: out <= 16'hFC79;    16'd28423: out <= 16'h0193;
    16'd28424: out <= 16'h042C;    16'd28425: out <= 16'hF95A;    16'd28426: out <= 16'h012A;    16'd28427: out <= 16'hFC7A;
    16'd28428: out <= 16'hFD2A;    16'd28429: out <= 16'h0A0B;    16'd28430: out <= 16'h01A7;    16'd28431: out <= 16'hFEE4;
    16'd28432: out <= 16'h041C;    16'd28433: out <= 16'hFDEA;    16'd28434: out <= 16'hFDEF;    16'd28435: out <= 16'h0702;
    16'd28436: out <= 16'h003B;    16'd28437: out <= 16'hFCDF;    16'd28438: out <= 16'h039E;    16'd28439: out <= 16'hFFA2;
    16'd28440: out <= 16'h01C8;    16'd28441: out <= 16'h0406;    16'd28442: out <= 16'h08BB;    16'd28443: out <= 16'h0385;
    16'd28444: out <= 16'h005D;    16'd28445: out <= 16'h0786;    16'd28446: out <= 16'hFBFB;    16'd28447: out <= 16'h0059;
    16'd28448: out <= 16'h0327;    16'd28449: out <= 16'h0357;    16'd28450: out <= 16'h09BF;    16'd28451: out <= 16'h03F3;
    16'd28452: out <= 16'hFD5D;    16'd28453: out <= 16'h0666;    16'd28454: out <= 16'h0742;    16'd28455: out <= 16'h0ABA;
    16'd28456: out <= 16'h09E8;    16'd28457: out <= 16'hFE72;    16'd28458: out <= 16'h07F3;    16'd28459: out <= 16'h0629;
    16'd28460: out <= 16'hFF4A;    16'd28461: out <= 16'hF8B2;    16'd28462: out <= 16'h0968;    16'd28463: out <= 16'h0340;
    16'd28464: out <= 16'h0058;    16'd28465: out <= 16'h033F;    16'd28466: out <= 16'h03FC;    16'd28467: out <= 16'h071F;
    16'd28468: out <= 16'h0E0C;    16'd28469: out <= 16'h0306;    16'd28470: out <= 16'h01B0;    16'd28471: out <= 16'h0269;
    16'd28472: out <= 16'h03D9;    16'd28473: out <= 16'h0170;    16'd28474: out <= 16'h0174;    16'd28475: out <= 16'h0065;
    16'd28476: out <= 16'h05F3;    16'd28477: out <= 16'h0AED;    16'd28478: out <= 16'h07CF;    16'd28479: out <= 16'h046D;
    16'd28480: out <= 16'h03A6;    16'd28481: out <= 16'h03F5;    16'd28482: out <= 16'h02E4;    16'd28483: out <= 16'hFFFD;
    16'd28484: out <= 16'hFFDB;    16'd28485: out <= 16'h081D;    16'd28486: out <= 16'h0528;    16'd28487: out <= 16'h04BB;
    16'd28488: out <= 16'h05C8;    16'd28489: out <= 16'h049A;    16'd28490: out <= 16'h0E4C;    16'd28491: out <= 16'h0175;
    16'd28492: out <= 16'h0085;    16'd28493: out <= 16'h0383;    16'd28494: out <= 16'h00F1;    16'd28495: out <= 16'h0418;
    16'd28496: out <= 16'h077A;    16'd28497: out <= 16'h0122;    16'd28498: out <= 16'h067C;    16'd28499: out <= 16'h02BC;
    16'd28500: out <= 16'h02DA;    16'd28501: out <= 16'h016D;    16'd28502: out <= 16'h0437;    16'd28503: out <= 16'h036C;
    16'd28504: out <= 16'h04A6;    16'd28505: out <= 16'h04D3;    16'd28506: out <= 16'hFD7A;    16'd28507: out <= 16'hFD95;
    16'd28508: out <= 16'h00A8;    16'd28509: out <= 16'h0581;    16'd28510: out <= 16'h04B8;    16'd28511: out <= 16'h022F;
    16'd28512: out <= 16'h01CC;    16'd28513: out <= 16'hFFC7;    16'd28514: out <= 16'h0181;    16'd28515: out <= 16'h04CD;
    16'd28516: out <= 16'h0313;    16'd28517: out <= 16'h0410;    16'd28518: out <= 16'h00A4;    16'd28519: out <= 16'h041B;
    16'd28520: out <= 16'hFFD9;    16'd28521: out <= 16'h03DE;    16'd28522: out <= 16'h05E1;    16'd28523: out <= 16'h09B5;
    16'd28524: out <= 16'h00E0;    16'd28525: out <= 16'h06FC;    16'd28526: out <= 16'h029C;    16'd28527: out <= 16'h0AF8;
    16'd28528: out <= 16'h0637;    16'd28529: out <= 16'h0525;    16'd28530: out <= 16'h06B2;    16'd28531: out <= 16'h01C3;
    16'd28532: out <= 16'h01CC;    16'd28533: out <= 16'h03A9;    16'd28534: out <= 16'h05A7;    16'd28535: out <= 16'h0414;
    16'd28536: out <= 16'h046F;    16'd28537: out <= 16'h0493;    16'd28538: out <= 16'h087F;    16'd28539: out <= 16'h08D4;
    16'd28540: out <= 16'h006C;    16'd28541: out <= 16'h020E;    16'd28542: out <= 16'h084D;    16'd28543: out <= 16'hFFF1;
    16'd28544: out <= 16'hFE18;    16'd28545: out <= 16'h02E8;    16'd28546: out <= 16'h00DA;    16'd28547: out <= 16'h051E;
    16'd28548: out <= 16'h03D7;    16'd28549: out <= 16'h022D;    16'd28550: out <= 16'h01B4;    16'd28551: out <= 16'h048C;
    16'd28552: out <= 16'h0854;    16'd28553: out <= 16'h053A;    16'd28554: out <= 16'h067B;    16'd28555: out <= 16'h08AA;
    16'd28556: out <= 16'h0302;    16'd28557: out <= 16'hFFF9;    16'd28558: out <= 16'h04F3;    16'd28559: out <= 16'h0457;
    16'd28560: out <= 16'h0478;    16'd28561: out <= 16'h0253;    16'd28562: out <= 16'h03A3;    16'd28563: out <= 16'h0FFE;
    16'd28564: out <= 16'h02D7;    16'd28565: out <= 16'h0060;    16'd28566: out <= 16'h030E;    16'd28567: out <= 16'h0433;
    16'd28568: out <= 16'hFDA5;    16'd28569: out <= 16'h06D7;    16'd28570: out <= 16'hFED0;    16'd28571: out <= 16'h022F;
    16'd28572: out <= 16'h084B;    16'd28573: out <= 16'hFE3C;    16'd28574: out <= 16'hFE52;    16'd28575: out <= 16'h018B;
    16'd28576: out <= 16'h07E0;    16'd28577: out <= 16'h0430;    16'd28578: out <= 16'h0748;    16'd28579: out <= 16'h0288;
    16'd28580: out <= 16'hFFA5;    16'd28581: out <= 16'h0391;    16'd28582: out <= 16'h05E1;    16'd28583: out <= 16'h05D3;
    16'd28584: out <= 16'h0C03;    16'd28585: out <= 16'h0B72;    16'd28586: out <= 16'h02D1;    16'd28587: out <= 16'h0E31;
    16'd28588: out <= 16'h0759;    16'd28589: out <= 16'h0094;    16'd28590: out <= 16'h07FD;    16'd28591: out <= 16'hFF63;
    16'd28592: out <= 16'hFF41;    16'd28593: out <= 16'h015E;    16'd28594: out <= 16'hFFEF;    16'd28595: out <= 16'h08D5;
    16'd28596: out <= 16'h0210;    16'd28597: out <= 16'hFE8D;    16'd28598: out <= 16'hFD5F;    16'd28599: out <= 16'h05C5;
    16'd28600: out <= 16'h0351;    16'd28601: out <= 16'h08D9;    16'd28602: out <= 16'h0332;    16'd28603: out <= 16'h04C5;
    16'd28604: out <= 16'hFE46;    16'd28605: out <= 16'h0A32;    16'd28606: out <= 16'h09CA;    16'd28607: out <= 16'hFCD5;
    16'd28608: out <= 16'hFF6B;    16'd28609: out <= 16'h09A5;    16'd28610: out <= 16'h0388;    16'd28611: out <= 16'h00DE;
    16'd28612: out <= 16'hFFF8;    16'd28613: out <= 16'h00DD;    16'd28614: out <= 16'h0092;    16'd28615: out <= 16'h003F;
    16'd28616: out <= 16'h0102;    16'd28617: out <= 16'h0AC4;    16'd28618: out <= 16'h00D3;    16'd28619: out <= 16'h04A0;
    16'd28620: out <= 16'h09A6;    16'd28621: out <= 16'h0777;    16'd28622: out <= 16'h0443;    16'd28623: out <= 16'h0085;
    16'd28624: out <= 16'h03D7;    16'd28625: out <= 16'hFE74;    16'd28626: out <= 16'hFFCA;    16'd28627: out <= 16'h065B;
    16'd28628: out <= 16'h0585;    16'd28629: out <= 16'h0500;    16'd28630: out <= 16'h0653;    16'd28631: out <= 16'h0393;
    16'd28632: out <= 16'h06ED;    16'd28633: out <= 16'hFF50;    16'd28634: out <= 16'hF2C7;    16'd28635: out <= 16'h0178;
    16'd28636: out <= 16'hFF54;    16'd28637: out <= 16'h024D;    16'd28638: out <= 16'h00F8;    16'd28639: out <= 16'h00D9;
    16'd28640: out <= 16'hFDBF;    16'd28641: out <= 16'h01DC;    16'd28642: out <= 16'hFEE3;    16'd28643: out <= 16'hFC91;
    16'd28644: out <= 16'hF755;    16'd28645: out <= 16'hFAF6;    16'd28646: out <= 16'hFDAE;    16'd28647: out <= 16'hF907;
    16'd28648: out <= 16'h0458;    16'd28649: out <= 16'hFAB4;    16'd28650: out <= 16'h0982;    16'd28651: out <= 16'hFE9F;
    16'd28652: out <= 16'h0369;    16'd28653: out <= 16'hFA4D;    16'd28654: out <= 16'h0388;    16'd28655: out <= 16'h0113;
    16'd28656: out <= 16'h00C5;    16'd28657: out <= 16'h024F;    16'd28658: out <= 16'h01B7;    16'd28659: out <= 16'hFEAC;
    16'd28660: out <= 16'h006D;    16'd28661: out <= 16'hF556;    16'd28662: out <= 16'h00FF;    16'd28663: out <= 16'hFFE5;
    16'd28664: out <= 16'h065C;    16'd28665: out <= 16'h03AF;    16'd28666: out <= 16'hFE0F;    16'd28667: out <= 16'hFE4F;
    16'd28668: out <= 16'hFF9D;    16'd28669: out <= 16'hFC4C;    16'd28670: out <= 16'h02EA;    16'd28671: out <= 16'hFF9B;
    16'd28672: out <= 16'h01EB;    16'd28673: out <= 16'h0131;    16'd28674: out <= 16'hFE9F;    16'd28675: out <= 16'hFA34;
    16'd28676: out <= 16'h040D;    16'd28677: out <= 16'hF875;    16'd28678: out <= 16'hFE16;    16'd28679: out <= 16'h04C9;
    16'd28680: out <= 16'hFB74;    16'd28681: out <= 16'h02C1;    16'd28682: out <= 16'h0051;    16'd28683: out <= 16'h001B;
    16'd28684: out <= 16'hFFF3;    16'd28685: out <= 16'h0179;    16'd28686: out <= 16'h02AC;    16'd28687: out <= 16'hF92C;
    16'd28688: out <= 16'h0383;    16'd28689: out <= 16'hFD37;    16'd28690: out <= 16'h08B2;    16'd28691: out <= 16'hFD0E;
    16'd28692: out <= 16'hFE7C;    16'd28693: out <= 16'hF7ED;    16'd28694: out <= 16'h018F;    16'd28695: out <= 16'hFEA7;
    16'd28696: out <= 16'h0533;    16'd28697: out <= 16'h018A;    16'd28698: out <= 16'h041F;    16'd28699: out <= 16'h012C;
    16'd28700: out <= 16'h05E4;    16'd28701: out <= 16'h071F;    16'd28702: out <= 16'hF97A;    16'd28703: out <= 16'h054B;
    16'd28704: out <= 16'h02DA;    16'd28705: out <= 16'h098A;    16'd28706: out <= 16'h06AD;    16'd28707: out <= 16'h0A1E;
    16'd28708: out <= 16'h0533;    16'd28709: out <= 16'hFFCF;    16'd28710: out <= 16'h08C1;    16'd28711: out <= 16'h0031;
    16'd28712: out <= 16'h0093;    16'd28713: out <= 16'h04DB;    16'd28714: out <= 16'h0594;    16'd28715: out <= 16'h0540;
    16'd28716: out <= 16'h04F9;    16'd28717: out <= 16'h049A;    16'd28718: out <= 16'h04C3;    16'd28719: out <= 16'h04C7;
    16'd28720: out <= 16'h07A8;    16'd28721: out <= 16'h00A3;    16'd28722: out <= 16'h0616;    16'd28723: out <= 16'h06D5;
    16'd28724: out <= 16'hFF83;    16'd28725: out <= 16'h0524;    16'd28726: out <= 16'hFF18;    16'd28727: out <= 16'h05CF;
    16'd28728: out <= 16'h0322;    16'd28729: out <= 16'hFF27;    16'd28730: out <= 16'h069D;    16'd28731: out <= 16'h0453;
    16'd28732: out <= 16'h0532;    16'd28733: out <= 16'h01CD;    16'd28734: out <= 16'h0167;    16'd28735: out <= 16'hFE14;
    16'd28736: out <= 16'h0054;    16'd28737: out <= 16'h0490;    16'd28738: out <= 16'hFE4C;    16'd28739: out <= 16'h0041;
    16'd28740: out <= 16'h038F;    16'd28741: out <= 16'h0890;    16'd28742: out <= 16'h06AF;    16'd28743: out <= 16'h049B;
    16'd28744: out <= 16'hFE94;    16'd28745: out <= 16'h01C1;    16'd28746: out <= 16'hFFBD;    16'd28747: out <= 16'h06F8;
    16'd28748: out <= 16'h03E4;    16'd28749: out <= 16'h08BD;    16'd28750: out <= 16'h040F;    16'd28751: out <= 16'h06D0;
    16'd28752: out <= 16'h0651;    16'd28753: out <= 16'h03C3;    16'd28754: out <= 16'h06D2;    16'd28755: out <= 16'h052A;
    16'd28756: out <= 16'h0733;    16'd28757: out <= 16'h0508;    16'd28758: out <= 16'h01E5;    16'd28759: out <= 16'h0258;
    16'd28760: out <= 16'h07E1;    16'd28761: out <= 16'h0225;    16'd28762: out <= 16'h0300;    16'd28763: out <= 16'h0236;
    16'd28764: out <= 16'hFEB4;    16'd28765: out <= 16'hFE22;    16'd28766: out <= 16'h088A;    16'd28767: out <= 16'h0E43;
    16'd28768: out <= 16'h062F;    16'd28769: out <= 16'h0134;    16'd28770: out <= 16'h05FD;    16'd28771: out <= 16'hFE2E;
    16'd28772: out <= 16'h0011;    16'd28773: out <= 16'h0A10;    16'd28774: out <= 16'h076E;    16'd28775: out <= 16'h03F5;
    16'd28776: out <= 16'h069C;    16'd28777: out <= 16'hFAAA;    16'd28778: out <= 16'h04FE;    16'd28779: out <= 16'h05AE;
    16'd28780: out <= 16'h04D6;    16'd28781: out <= 16'h0495;    16'd28782: out <= 16'h0859;    16'd28783: out <= 16'h0297;
    16'd28784: out <= 16'hFE4C;    16'd28785: out <= 16'h0163;    16'd28786: out <= 16'h01DA;    16'd28787: out <= 16'h04E3;
    16'd28788: out <= 16'h0368;    16'd28789: out <= 16'h0338;    16'd28790: out <= 16'h058E;    16'd28791: out <= 16'h03A4;
    16'd28792: out <= 16'h053A;    16'd28793: out <= 16'h05CC;    16'd28794: out <= 16'h0171;    16'd28795: out <= 16'h0856;
    16'd28796: out <= 16'h0843;    16'd28797: out <= 16'h02AF;    16'd28798: out <= 16'hFE61;    16'd28799: out <= 16'h01C7;
    16'd28800: out <= 16'h04E8;    16'd28801: out <= 16'h051F;    16'd28802: out <= 16'h0096;    16'd28803: out <= 16'hFDBA;
    16'd28804: out <= 16'h006A;    16'd28805: out <= 16'h02D7;    16'd28806: out <= 16'h0540;    16'd28807: out <= 16'h0476;
    16'd28808: out <= 16'h02B7;    16'd28809: out <= 16'h02FA;    16'd28810: out <= 16'h068C;    16'd28811: out <= 16'h038B;
    16'd28812: out <= 16'hFF02;    16'd28813: out <= 16'h01BD;    16'd28814: out <= 16'h079A;    16'd28815: out <= 16'hFF3C;
    16'd28816: out <= 16'h0026;    16'd28817: out <= 16'h03A6;    16'd28818: out <= 16'hF77A;    16'd28819: out <= 16'h008C;
    16'd28820: out <= 16'h0551;    16'd28821: out <= 16'h0754;    16'd28822: out <= 16'h04F3;    16'd28823: out <= 16'h0358;
    16'd28824: out <= 16'h00FD;    16'd28825: out <= 16'h03CF;    16'd28826: out <= 16'h0545;    16'd28827: out <= 16'h0331;
    16'd28828: out <= 16'h05B7;    16'd28829: out <= 16'hFFF8;    16'd28830: out <= 16'h0AD4;    16'd28831: out <= 16'h0CB5;
    16'd28832: out <= 16'hFE52;    16'd28833: out <= 16'hFFBB;    16'd28834: out <= 16'hFE1B;    16'd28835: out <= 16'h0233;
    16'd28836: out <= 16'h03A4;    16'd28837: out <= 16'h03A6;    16'd28838: out <= 16'h0069;    16'd28839: out <= 16'h001C;
    16'd28840: out <= 16'hFC84;    16'd28841: out <= 16'h0435;    16'd28842: out <= 16'h0140;    16'd28843: out <= 16'h00F3;
    16'd28844: out <= 16'h06BE;    16'd28845: out <= 16'h0263;    16'd28846: out <= 16'h01BD;    16'd28847: out <= 16'h0948;
    16'd28848: out <= 16'hFE03;    16'd28849: out <= 16'h0162;    16'd28850: out <= 16'h0105;    16'd28851: out <= 16'h0473;
    16'd28852: out <= 16'h0451;    16'd28853: out <= 16'h059A;    16'd28854: out <= 16'h03F1;    16'd28855: out <= 16'h03F3;
    16'd28856: out <= 16'h066D;    16'd28857: out <= 16'h02AE;    16'd28858: out <= 16'h081E;    16'd28859: out <= 16'h0305;
    16'd28860: out <= 16'h018B;    16'd28861: out <= 16'h04A1;    16'd28862: out <= 16'h06A7;    16'd28863: out <= 16'h02BC;
    16'd28864: out <= 16'h009D;    16'd28865: out <= 16'h01B0;    16'd28866: out <= 16'hFE72;    16'd28867: out <= 16'h0BB2;
    16'd28868: out <= 16'h0873;    16'd28869: out <= 16'hFB9D;    16'd28870: out <= 16'h07C1;    16'd28871: out <= 16'h0101;
    16'd28872: out <= 16'h00FF;    16'd28873: out <= 16'h026D;    16'd28874: out <= 16'h035B;    16'd28875: out <= 16'h067C;
    16'd28876: out <= 16'h0889;    16'd28877: out <= 16'h0091;    16'd28878: out <= 16'hF9F5;    16'd28879: out <= 16'h0080;
    16'd28880: out <= 16'hFFE9;    16'd28881: out <= 16'h0311;    16'd28882: out <= 16'h03F6;    16'd28883: out <= 16'h017A;
    16'd28884: out <= 16'h0C5D;    16'd28885: out <= 16'h04D9;    16'd28886: out <= 16'h0152;    16'd28887: out <= 16'h05FC;
    16'd28888: out <= 16'h03C1;    16'd28889: out <= 16'hFEF2;    16'd28890: out <= 16'hFD93;    16'd28891: out <= 16'hFF9C;
    16'd28892: out <= 16'hFB21;    16'd28893: out <= 16'h0428;    16'd28894: out <= 16'hF89B;    16'd28895: out <= 16'h0300;
    16'd28896: out <= 16'h0912;    16'd28897: out <= 16'h0196;    16'd28898: out <= 16'hFE09;    16'd28899: out <= 16'h0262;
    16'd28900: out <= 16'h02A1;    16'd28901: out <= 16'h05FF;    16'd28902: out <= 16'hFE04;    16'd28903: out <= 16'h0087;
    16'd28904: out <= 16'h007B;    16'd28905: out <= 16'hF964;    16'd28906: out <= 16'hFF76;    16'd28907: out <= 16'hFDF6;
    16'd28908: out <= 16'h0253;    16'd28909: out <= 16'hFFAF;    16'd28910: out <= 16'h08A2;    16'd28911: out <= 16'hFDAA;
    16'd28912: out <= 16'h048D;    16'd28913: out <= 16'hFF15;    16'd28914: out <= 16'h047D;    16'd28915: out <= 16'h00A7;
    16'd28916: out <= 16'h08CC;    16'd28917: out <= 16'hFC94;    16'd28918: out <= 16'h0244;    16'd28919: out <= 16'h0874;
    16'd28920: out <= 16'hFC85;    16'd28921: out <= 16'hFB6C;    16'd28922: out <= 16'h026D;    16'd28923: out <= 16'h009B;
    16'd28924: out <= 16'hFD02;    16'd28925: out <= 16'hFE1A;    16'd28926: out <= 16'hFB45;    16'd28927: out <= 16'h02B0;
    16'd28928: out <= 16'h05DB;    16'd28929: out <= 16'h0432;    16'd28930: out <= 16'h006B;    16'd28931: out <= 16'hFEFE;
    16'd28932: out <= 16'h0127;    16'd28933: out <= 16'hFE87;    16'd28934: out <= 16'hFFB5;    16'd28935: out <= 16'hFDE9;
    16'd28936: out <= 16'h0557;    16'd28937: out <= 16'h0183;    16'd28938: out <= 16'hF5AE;    16'd28939: out <= 16'hFB9E;
    16'd28940: out <= 16'hFA4F;    16'd28941: out <= 16'h050C;    16'd28942: out <= 16'hFCDE;    16'd28943: out <= 16'hFAB8;
    16'd28944: out <= 16'h02F5;    16'd28945: out <= 16'h009A;    16'd28946: out <= 16'h00C9;    16'd28947: out <= 16'hFE95;
    16'd28948: out <= 16'hF936;    16'd28949: out <= 16'h01BA;    16'd28950: out <= 16'h011B;    16'd28951: out <= 16'h068D;
    16'd28952: out <= 16'h0598;    16'd28953: out <= 16'h048C;    16'd28954: out <= 16'h00B1;    16'd28955: out <= 16'h0452;
    16'd28956: out <= 16'h057B;    16'd28957: out <= 16'h084A;    16'd28958: out <= 16'h0215;    16'd28959: out <= 16'h01DE;
    16'd28960: out <= 16'h00F0;    16'd28961: out <= 16'h088F;    16'd28962: out <= 16'h002D;    16'd28963: out <= 16'h0406;
    16'd28964: out <= 16'h04AB;    16'd28965: out <= 16'h0258;    16'd28966: out <= 16'h0298;    16'd28967: out <= 16'h0311;
    16'd28968: out <= 16'h0783;    16'd28969: out <= 16'h0594;    16'd28970: out <= 16'h0505;    16'd28971: out <= 16'h0A16;
    16'd28972: out <= 16'hFCC5;    16'd28973: out <= 16'h07D3;    16'd28974: out <= 16'h0799;    16'd28975: out <= 16'h01A6;
    16'd28976: out <= 16'h03C7;    16'd28977: out <= 16'h00D1;    16'd28978: out <= 16'h02AE;    16'd28979: out <= 16'h061A;
    16'd28980: out <= 16'hFC9E;    16'd28981: out <= 16'h05C3;    16'd28982: out <= 16'h073A;    16'd28983: out <= 16'h017E;
    16'd28984: out <= 16'h0690;    16'd28985: out <= 16'h074E;    16'd28986: out <= 16'h013F;    16'd28987: out <= 16'h11B3;
    16'd28988: out <= 16'h083E;    16'd28989: out <= 16'hFF88;    16'd28990: out <= 16'hFE91;    16'd28991: out <= 16'h072C;
    16'd28992: out <= 16'h04FB;    16'd28993: out <= 16'h027A;    16'd28994: out <= 16'hFDB9;    16'd28995: out <= 16'hFFFA;
    16'd28996: out <= 16'h0593;    16'd28997: out <= 16'h0509;    16'd28998: out <= 16'h04F0;    16'd28999: out <= 16'h0549;
    16'd29000: out <= 16'h0656;    16'd29001: out <= 16'h0807;    16'd29002: out <= 16'h00B0;    16'd29003: out <= 16'hFC50;
    16'd29004: out <= 16'h0082;    16'd29005: out <= 16'h0504;    16'd29006: out <= 16'h06A1;    16'd29007: out <= 16'h0DB3;
    16'd29008: out <= 16'h0282;    16'd29009: out <= 16'h07B6;    16'd29010: out <= 16'h048F;    16'd29011: out <= 16'h0AF3;
    16'd29012: out <= 16'h0117;    16'd29013: out <= 16'h0057;    16'd29014: out <= 16'h0137;    16'd29015: out <= 16'h0911;
    16'd29016: out <= 16'h09EA;    16'd29017: out <= 16'h03BD;    16'd29018: out <= 16'h04D0;    16'd29019: out <= 16'hFDB4;
    16'd29020: out <= 16'hFD8C;    16'd29021: out <= 16'hFF6A;    16'd29022: out <= 16'h0AE3;    16'd29023: out <= 16'h0153;
    16'd29024: out <= 16'h0657;    16'd29025: out <= 16'h0B03;    16'd29026: out <= 16'hFFDB;    16'd29027: out <= 16'h069E;
    16'd29028: out <= 16'h01B5;    16'd29029: out <= 16'h0495;    16'd29030: out <= 16'h04D8;    16'd29031: out <= 16'h059B;
    16'd29032: out <= 16'h045B;    16'd29033: out <= 16'hFB21;    16'd29034: out <= 16'h0B7C;    16'd29035: out <= 16'h0C6F;
    16'd29036: out <= 16'hFF6C;    16'd29037: out <= 16'h00EA;    16'd29038: out <= 16'h04BD;    16'd29039: out <= 16'h0532;
    16'd29040: out <= 16'h086B;    16'd29041: out <= 16'h036B;    16'd29042: out <= 16'hFD9E;    16'd29043: out <= 16'h02D7;
    16'd29044: out <= 16'hFF13;    16'd29045: out <= 16'h07FD;    16'd29046: out <= 16'h04BB;    16'd29047: out <= 16'h0A95;
    16'd29048: out <= 16'h04B2;    16'd29049: out <= 16'h035A;    16'd29050: out <= 16'h0276;    16'd29051: out <= 16'hFC2D;
    16'd29052: out <= 16'h0350;    16'd29053: out <= 16'h0837;    16'd29054: out <= 16'h0487;    16'd29055: out <= 16'h0795;
    16'd29056: out <= 16'h02C5;    16'd29057: out <= 16'hF9A4;    16'd29058: out <= 16'h01E4;    16'd29059: out <= 16'h0431;
    16'd29060: out <= 16'h0399;    16'd29061: out <= 16'h031B;    16'd29062: out <= 16'hFAAE;    16'd29063: out <= 16'h04E7;
    16'd29064: out <= 16'hFDD6;    16'd29065: out <= 16'h00CE;    16'd29066: out <= 16'h04B0;    16'd29067: out <= 16'h041D;
    16'd29068: out <= 16'h08A6;    16'd29069: out <= 16'h063A;    16'd29070: out <= 16'h057A;    16'd29071: out <= 16'h019A;
    16'd29072: out <= 16'h03B5;    16'd29073: out <= 16'h0264;    16'd29074: out <= 16'h0214;    16'd29075: out <= 16'hFEB5;
    16'd29076: out <= 16'h059C;    16'd29077: out <= 16'h0BFA;    16'd29078: out <= 16'h0409;    16'd29079: out <= 16'h0417;
    16'd29080: out <= 16'h053B;    16'd29081: out <= 16'h06D0;    16'd29082: out <= 16'h00A4;    16'd29083: out <= 16'h0083;
    16'd29084: out <= 16'hFF34;    16'd29085: out <= 16'hFD3F;    16'd29086: out <= 16'h024E;    16'd29087: out <= 16'h0286;
    16'd29088: out <= 16'h00AD;    16'd29089: out <= 16'h05F1;    16'd29090: out <= 16'hFF9F;    16'd29091: out <= 16'h0631;
    16'd29092: out <= 16'h03EE;    16'd29093: out <= 16'h0226;    16'd29094: out <= 16'hFF1F;    16'd29095: out <= 16'h041E;
    16'd29096: out <= 16'h02DF;    16'd29097: out <= 16'h0500;    16'd29098: out <= 16'h0684;    16'd29099: out <= 16'h035E;
    16'd29100: out <= 16'h0653;    16'd29101: out <= 16'h0494;    16'd29102: out <= 16'h088D;    16'd29103: out <= 16'hFCD1;
    16'd29104: out <= 16'h0299;    16'd29105: out <= 16'hFAE5;    16'd29106: out <= 16'hFECD;    16'd29107: out <= 16'h0314;
    16'd29108: out <= 16'h0373;    16'd29109: out <= 16'hFCB9;    16'd29110: out <= 16'h0184;    16'd29111: out <= 16'h0572;
    16'd29112: out <= 16'h0862;    16'd29113: out <= 16'hF7D0;    16'd29114: out <= 16'h0515;    16'd29115: out <= 16'h00E0;
    16'd29116: out <= 16'h042D;    16'd29117: out <= 16'hFED9;    16'd29118: out <= 16'h03A8;    16'd29119: out <= 16'hFD8F;
    16'd29120: out <= 16'h01A1;    16'd29121: out <= 16'h016F;    16'd29122: out <= 16'h045A;    16'd29123: out <= 16'h0750;
    16'd29124: out <= 16'h0336;    16'd29125: out <= 16'hFF90;    16'd29126: out <= 16'h0823;    16'd29127: out <= 16'hFD7D;
    16'd29128: out <= 16'h00B1;    16'd29129: out <= 16'h08C9;    16'd29130: out <= 16'h038B;    16'd29131: out <= 16'h07B4;
    16'd29132: out <= 16'h04D3;    16'd29133: out <= 16'h0316;    16'd29134: out <= 16'h0499;    16'd29135: out <= 16'h0484;
    16'd29136: out <= 16'h0207;    16'd29137: out <= 16'hFB96;    16'd29138: out <= 16'h03AB;    16'd29139: out <= 16'h0A62;
    16'd29140: out <= 16'h035E;    16'd29141: out <= 16'hFAE2;    16'd29142: out <= 16'h02C8;    16'd29143: out <= 16'h0797;
    16'd29144: out <= 16'h0AAC;    16'd29145: out <= 16'h026E;    16'd29146: out <= 16'h030B;    16'd29147: out <= 16'h0288;
    16'd29148: out <= 16'hFAE9;    16'd29149: out <= 16'h0391;    16'd29150: out <= 16'h0420;    16'd29151: out <= 16'h005B;
    16'd29152: out <= 16'h0188;    16'd29153: out <= 16'hFD58;    16'd29154: out <= 16'hF817;    16'd29155: out <= 16'hFBF5;
    16'd29156: out <= 16'hFE05;    16'd29157: out <= 16'hFE15;    16'd29158: out <= 16'hFD36;    16'd29159: out <= 16'h00D3;
    16'd29160: out <= 16'hFD0B;    16'd29161: out <= 16'hFD2A;    16'd29162: out <= 16'hFB68;    16'd29163: out <= 16'hFF35;
    16'd29164: out <= 16'hFD58;    16'd29165: out <= 16'hF956;    16'd29166: out <= 16'h03FA;    16'd29167: out <= 16'h005B;
    16'd29168: out <= 16'h0624;    16'd29169: out <= 16'h00FF;    16'd29170: out <= 16'h086C;    16'd29171: out <= 16'hFECE;
    16'd29172: out <= 16'h0684;    16'd29173: out <= 16'hFC1E;    16'd29174: out <= 16'h05A8;    16'd29175: out <= 16'hFD8B;
    16'd29176: out <= 16'hFFD9;    16'd29177: out <= 16'h0023;    16'd29178: out <= 16'hF7A0;    16'd29179: out <= 16'h04DC;
    16'd29180: out <= 16'h05C7;    16'd29181: out <= 16'hF703;    16'd29182: out <= 16'h013D;    16'd29183: out <= 16'h0049;
    16'd29184: out <= 16'hFC0F;    16'd29185: out <= 16'h062F;    16'd29186: out <= 16'h0657;    16'd29187: out <= 16'h037A;
    16'd29188: out <= 16'hFC0B;    16'd29189: out <= 16'hFE2F;    16'd29190: out <= 16'h03FF;    16'd29191: out <= 16'h0511;
    16'd29192: out <= 16'h01EC;    16'd29193: out <= 16'hF77F;    16'd29194: out <= 16'h0042;    16'd29195: out <= 16'h0285;
    16'd29196: out <= 16'hFBBD;    16'd29197: out <= 16'hF8F3;    16'd29198: out <= 16'h03A0;    16'd29199: out <= 16'h0284;
    16'd29200: out <= 16'h00C6;    16'd29201: out <= 16'hFDA9;    16'd29202: out <= 16'hFF78;    16'd29203: out <= 16'hFBA6;
    16'd29204: out <= 16'hFC0E;    16'd29205: out <= 16'hFEDA;    16'd29206: out <= 16'h0714;    16'd29207: out <= 16'h0027;
    16'd29208: out <= 16'hFE59;    16'd29209: out <= 16'h0E75;    16'd29210: out <= 16'h0479;    16'd29211: out <= 16'h080B;
    16'd29212: out <= 16'h08F5;    16'd29213: out <= 16'h03A3;    16'd29214: out <= 16'h0998;    16'd29215: out <= 16'hFD58;
    16'd29216: out <= 16'h018D;    16'd29217: out <= 16'h0536;    16'd29218: out <= 16'h02E2;    16'd29219: out <= 16'h0626;
    16'd29220: out <= 16'h05DB;    16'd29221: out <= 16'h0749;    16'd29222: out <= 16'hFBC9;    16'd29223: out <= 16'h0588;
    16'd29224: out <= 16'h00D5;    16'd29225: out <= 16'hFD6D;    16'd29226: out <= 16'h03A3;    16'd29227: out <= 16'h0475;
    16'd29228: out <= 16'h017C;    16'd29229: out <= 16'h0AB8;    16'd29230: out <= 16'h03AF;    16'd29231: out <= 16'h0950;
    16'd29232: out <= 16'h0682;    16'd29233: out <= 16'h0239;    16'd29234: out <= 16'h0A31;    16'd29235: out <= 16'h056C;
    16'd29236: out <= 16'hFFD4;    16'd29237: out <= 16'h0101;    16'd29238: out <= 16'h0463;    16'd29239: out <= 16'h005C;
    16'd29240: out <= 16'h02EA;    16'd29241: out <= 16'hFE9E;    16'd29242: out <= 16'h0328;    16'd29243: out <= 16'h032B;
    16'd29244: out <= 16'h00A6;    16'd29245: out <= 16'hFFA7;    16'd29246: out <= 16'h05ED;    16'd29247: out <= 16'h039E;
    16'd29248: out <= 16'hFFF3;    16'd29249: out <= 16'hFED3;    16'd29250: out <= 16'h083B;    16'd29251: out <= 16'h0231;
    16'd29252: out <= 16'h04BD;    16'd29253: out <= 16'h086E;    16'd29254: out <= 16'hFCC8;    16'd29255: out <= 16'hFFE5;
    16'd29256: out <= 16'hFD96;    16'd29257: out <= 16'h0509;    16'd29258: out <= 16'h05DB;    16'd29259: out <= 16'hFFDC;
    16'd29260: out <= 16'h03AD;    16'd29261: out <= 16'h04CC;    16'd29262: out <= 16'h095C;    16'd29263: out <= 16'h06B8;
    16'd29264: out <= 16'h04D8;    16'd29265: out <= 16'h05FC;    16'd29266: out <= 16'h0904;    16'd29267: out <= 16'h06BD;
    16'd29268: out <= 16'h04CA;    16'd29269: out <= 16'hFD53;    16'd29270: out <= 16'h066A;    16'd29271: out <= 16'h0707;
    16'd29272: out <= 16'h03D0;    16'd29273: out <= 16'hF7A3;    16'd29274: out <= 16'h0106;    16'd29275: out <= 16'h0077;
    16'd29276: out <= 16'h0811;    16'd29277: out <= 16'h08B8;    16'd29278: out <= 16'h0376;    16'd29279: out <= 16'h00B6;
    16'd29280: out <= 16'h04DD;    16'd29281: out <= 16'hFD45;    16'd29282: out <= 16'h074A;    16'd29283: out <= 16'h07B4;
    16'd29284: out <= 16'h02F6;    16'd29285: out <= 16'h0CD8;    16'd29286: out <= 16'h0186;    16'd29287: out <= 16'hFEA8;
    16'd29288: out <= 16'h0360;    16'd29289: out <= 16'h06DE;    16'd29290: out <= 16'hFD66;    16'd29291: out <= 16'h0330;
    16'd29292: out <= 16'h016F;    16'd29293: out <= 16'h0029;    16'd29294: out <= 16'h05DA;    16'd29295: out <= 16'h0363;
    16'd29296: out <= 16'hFCC9;    16'd29297: out <= 16'h0482;    16'd29298: out <= 16'h0494;    16'd29299: out <= 16'h03B5;
    16'd29300: out <= 16'h0D52;    16'd29301: out <= 16'h05C1;    16'd29302: out <= 16'hFF43;    16'd29303: out <= 16'h0581;
    16'd29304: out <= 16'h0539;    16'd29305: out <= 16'h050F;    16'd29306: out <= 16'h116C;    16'd29307: out <= 16'h02AB;
    16'd29308: out <= 16'h0304;    16'd29309: out <= 16'h0BC0;    16'd29310: out <= 16'h0120;    16'd29311: out <= 16'h0695;
    16'd29312: out <= 16'hF8F5;    16'd29313: out <= 16'h08C5;    16'd29314: out <= 16'h0073;    16'd29315: out <= 16'hFEFE;
    16'd29316: out <= 16'h0664;    16'd29317: out <= 16'h008B;    16'd29318: out <= 16'h0519;    16'd29319: out <= 16'hFF1F;
    16'd29320: out <= 16'h02DA;    16'd29321: out <= 16'h048C;    16'd29322: out <= 16'h07A0;    16'd29323: out <= 16'hFDBC;
    16'd29324: out <= 16'h0283;    16'd29325: out <= 16'h02C4;    16'd29326: out <= 16'h06F6;    16'd29327: out <= 16'h037E;
    16'd29328: out <= 16'h0372;    16'd29329: out <= 16'hFEC2;    16'd29330: out <= 16'h016E;    16'd29331: out <= 16'h02BE;
    16'd29332: out <= 16'hFF58;    16'd29333: out <= 16'h0729;    16'd29334: out <= 16'hFFA9;    16'd29335: out <= 16'h0148;
    16'd29336: out <= 16'h0277;    16'd29337: out <= 16'h0752;    16'd29338: out <= 16'h0865;    16'd29339: out <= 16'h0695;
    16'd29340: out <= 16'h0617;    16'd29341: out <= 16'h0548;    16'd29342: out <= 16'h03F5;    16'd29343: out <= 16'h0850;
    16'd29344: out <= 16'h027F;    16'd29345: out <= 16'hFE30;    16'd29346: out <= 16'h0392;    16'd29347: out <= 16'hFF63;
    16'd29348: out <= 16'h005B;    16'd29349: out <= 16'h02C4;    16'd29350: out <= 16'h04E4;    16'd29351: out <= 16'h02DD;
    16'd29352: out <= 16'h0033;    16'd29353: out <= 16'h0636;    16'd29354: out <= 16'h0911;    16'd29355: out <= 16'h0144;
    16'd29356: out <= 16'h0FD4;    16'd29357: out <= 16'h0872;    16'd29358: out <= 16'h064F;    16'd29359: out <= 16'h0173;
    16'd29360: out <= 16'hFE7C;    16'd29361: out <= 16'h02F2;    16'd29362: out <= 16'h0495;    16'd29363: out <= 16'h0C21;
    16'd29364: out <= 16'h02D9;    16'd29365: out <= 16'h085E;    16'd29366: out <= 16'hFFFA;    16'd29367: out <= 16'h0484;
    16'd29368: out <= 16'h02E9;    16'd29369: out <= 16'h04EF;    16'd29370: out <= 16'h0915;    16'd29371: out <= 16'h0582;
    16'd29372: out <= 16'h01AA;    16'd29373: out <= 16'h025A;    16'd29374: out <= 16'h0255;    16'd29375: out <= 16'h0447;
    16'd29376: out <= 16'h02DF;    16'd29377: out <= 16'h0AC3;    16'd29378: out <= 16'h0337;    16'd29379: out <= 16'h036B;
    16'd29380: out <= 16'h0465;    16'd29381: out <= 16'h0641;    16'd29382: out <= 16'h03E0;    16'd29383: out <= 16'h06D5;
    16'd29384: out <= 16'h01A9;    16'd29385: out <= 16'h0A51;    16'd29386: out <= 16'h0436;    16'd29387: out <= 16'hFFA8;
    16'd29388: out <= 16'h04FA;    16'd29389: out <= 16'h0120;    16'd29390: out <= 16'hFFC4;    16'd29391: out <= 16'h03AD;
    16'd29392: out <= 16'h076F;    16'd29393: out <= 16'h00DE;    16'd29394: out <= 16'h0625;    16'd29395: out <= 16'h035F;
    16'd29396: out <= 16'h0900;    16'd29397: out <= 16'h0A85;    16'd29398: out <= 16'hFFFC;    16'd29399: out <= 16'hFE59;
    16'd29400: out <= 16'h01D6;    16'd29401: out <= 16'h0572;    16'd29402: out <= 16'h0096;    16'd29403: out <= 16'hFC8A;
    16'd29404: out <= 16'hFF5D;    16'd29405: out <= 16'hFDD7;    16'd29406: out <= 16'hF83A;    16'd29407: out <= 16'h0016;
    16'd29408: out <= 16'h00DA;    16'd29409: out <= 16'hFFC5;    16'd29410: out <= 16'h00D5;    16'd29411: out <= 16'hF87E;
    16'd29412: out <= 16'hFE83;    16'd29413: out <= 16'hFC95;    16'd29414: out <= 16'hFDAC;    16'd29415: out <= 16'hFFAC;
    16'd29416: out <= 16'hFEB8;    16'd29417: out <= 16'h00B0;    16'd29418: out <= 16'hFA11;    16'd29419: out <= 16'h008E;
    16'd29420: out <= 16'hFD91;    16'd29421: out <= 16'hFC77;    16'd29422: out <= 16'h0486;    16'd29423: out <= 16'h069A;
    16'd29424: out <= 16'h05B8;    16'd29425: out <= 16'h0000;    16'd29426: out <= 16'h00AA;    16'd29427: out <= 16'hFA3B;
    16'd29428: out <= 16'h050B;    16'd29429: out <= 16'h049F;    16'd29430: out <= 16'h0138;    16'd29431: out <= 16'h0299;
    16'd29432: out <= 16'hFED3;    16'd29433: out <= 16'h0878;    16'd29434: out <= 16'hFEC5;    16'd29435: out <= 16'hF9A8;
    16'd29436: out <= 16'hFD65;    16'd29437: out <= 16'h0019;    16'd29438: out <= 16'hFC99;    16'd29439: out <= 16'hFC22;
    16'd29440: out <= 16'h052A;    16'd29441: out <= 16'h0035;    16'd29442: out <= 16'h02DE;    16'd29443: out <= 16'h0547;
    16'd29444: out <= 16'hF6F0;    16'd29445: out <= 16'h027D;    16'd29446: out <= 16'h0421;    16'd29447: out <= 16'h0095;
    16'd29448: out <= 16'hFAC5;    16'd29449: out <= 16'hF72C;    16'd29450: out <= 16'hFDCA;    16'd29451: out <= 16'hFB10;
    16'd29452: out <= 16'h0650;    16'd29453: out <= 16'hF9B2;    16'd29454: out <= 16'h06C5;    16'd29455: out <= 16'hFD0A;
    16'd29456: out <= 16'hFD57;    16'd29457: out <= 16'hFF18;    16'd29458: out <= 16'hFC33;    16'd29459: out <= 16'hFEC0;
    16'd29460: out <= 16'hFF62;    16'd29461: out <= 16'h09C8;    16'd29462: out <= 16'hFF63;    16'd29463: out <= 16'hFD0A;
    16'd29464: out <= 16'h02BF;    16'd29465: out <= 16'hFFA4;    16'd29466: out <= 16'h00C3;    16'd29467: out <= 16'h0559;
    16'd29468: out <= 16'h0B1D;    16'd29469: out <= 16'h047A;    16'd29470: out <= 16'h07E7;    16'd29471: out <= 16'hFF04;
    16'd29472: out <= 16'h06A4;    16'd29473: out <= 16'hFF94;    16'd29474: out <= 16'h04B5;    16'd29475: out <= 16'h0515;
    16'd29476: out <= 16'h0380;    16'd29477: out <= 16'hFF10;    16'd29478: out <= 16'h0BFB;    16'd29479: out <= 16'h073E;
    16'd29480: out <= 16'h0540;    16'd29481: out <= 16'h0E95;    16'd29482: out <= 16'h0340;    16'd29483: out <= 16'h00C5;
    16'd29484: out <= 16'hFDEF;    16'd29485: out <= 16'h03F9;    16'd29486: out <= 16'h020D;    16'd29487: out <= 16'h04DD;
    16'd29488: out <= 16'h0206;    16'd29489: out <= 16'h00AB;    16'd29490: out <= 16'h000C;    16'd29491: out <= 16'h007F;
    16'd29492: out <= 16'h0805;    16'd29493: out <= 16'h001E;    16'd29494: out <= 16'h0388;    16'd29495: out <= 16'h07AD;
    16'd29496: out <= 16'h06F5;    16'd29497: out <= 16'h0163;    16'd29498: out <= 16'h06C1;    16'd29499: out <= 16'h05D6;
    16'd29500: out <= 16'h0269;    16'd29501: out <= 16'h088A;    16'd29502: out <= 16'h075A;    16'd29503: out <= 16'h057B;
    16'd29504: out <= 16'h04E2;    16'd29505: out <= 16'h04BF;    16'd29506: out <= 16'h0680;    16'd29507: out <= 16'h0AC8;
    16'd29508: out <= 16'h01E1;    16'd29509: out <= 16'h0004;    16'd29510: out <= 16'h0508;    16'd29511: out <= 16'h0289;
    16'd29512: out <= 16'h03B1;    16'd29513: out <= 16'h017F;    16'd29514: out <= 16'h0784;    16'd29515: out <= 16'h0121;
    16'd29516: out <= 16'h01D4;    16'd29517: out <= 16'h053C;    16'd29518: out <= 16'h03B0;    16'd29519: out <= 16'h07AC;
    16'd29520: out <= 16'h0396;    16'd29521: out <= 16'h06A8;    16'd29522: out <= 16'h052D;    16'd29523: out <= 16'h04E6;
    16'd29524: out <= 16'h033A;    16'd29525: out <= 16'h0AAC;    16'd29526: out <= 16'h002B;    16'd29527: out <= 16'h027D;
    16'd29528: out <= 16'h0449;    16'd29529: out <= 16'h056B;    16'd29530: out <= 16'h0643;    16'd29531: out <= 16'h0335;
    16'd29532: out <= 16'h047C;    16'd29533: out <= 16'h0050;    16'd29534: out <= 16'h018D;    16'd29535: out <= 16'h07EF;
    16'd29536: out <= 16'h01A9;    16'd29537: out <= 16'h0215;    16'd29538: out <= 16'hFD7B;    16'd29539: out <= 16'h078A;
    16'd29540: out <= 16'h0624;    16'd29541: out <= 16'h0723;    16'd29542: out <= 16'h057B;    16'd29543: out <= 16'hFD6E;
    16'd29544: out <= 16'h0347;    16'd29545: out <= 16'h08B3;    16'd29546: out <= 16'h0556;    16'd29547: out <= 16'h0392;
    16'd29548: out <= 16'h0594;    16'd29549: out <= 16'h09BC;    16'd29550: out <= 16'h0670;    16'd29551: out <= 16'h0268;
    16'd29552: out <= 16'h03A3;    16'd29553: out <= 16'h099C;    16'd29554: out <= 16'h0381;    16'd29555: out <= 16'hFEEA;
    16'd29556: out <= 16'h0789;    16'd29557: out <= 16'h031D;    16'd29558: out <= 16'h01C8;    16'd29559: out <= 16'h03A9;
    16'd29560: out <= 16'hFE88;    16'd29561: out <= 16'h0BAF;    16'd29562: out <= 16'h03B0;    16'd29563: out <= 16'h043D;
    16'd29564: out <= 16'h0756;    16'd29565: out <= 16'h06EA;    16'd29566: out <= 16'h0209;    16'd29567: out <= 16'h0A36;
    16'd29568: out <= 16'h0951;    16'd29569: out <= 16'h0297;    16'd29570: out <= 16'h0251;    16'd29571: out <= 16'h09F1;
    16'd29572: out <= 16'h02B6;    16'd29573: out <= 16'h08D2;    16'd29574: out <= 16'h0822;    16'd29575: out <= 16'hFFA1;
    16'd29576: out <= 16'hFF84;    16'd29577: out <= 16'hFEB9;    16'd29578: out <= 16'h083F;    16'd29579: out <= 16'h0843;
    16'd29580: out <= 16'h0282;    16'd29581: out <= 16'h0467;    16'd29582: out <= 16'h048D;    16'd29583: out <= 16'h01C1;
    16'd29584: out <= 16'h07BC;    16'd29585: out <= 16'h00A0;    16'd29586: out <= 16'h0696;    16'd29587: out <= 16'h05D9;
    16'd29588: out <= 16'h07D2;    16'd29589: out <= 16'h0175;    16'd29590: out <= 16'hFF37;    16'd29591: out <= 16'h08B8;
    16'd29592: out <= 16'h0502;    16'd29593: out <= 16'h0875;    16'd29594: out <= 16'h03CC;    16'd29595: out <= 16'h07E6;
    16'd29596: out <= 16'hFEBB;    16'd29597: out <= 16'h02CB;    16'd29598: out <= 16'h037B;    16'd29599: out <= 16'h002A;
    16'd29600: out <= 16'h05C5;    16'd29601: out <= 16'h057E;    16'd29602: out <= 16'h02F0;    16'd29603: out <= 16'h04A8;
    16'd29604: out <= 16'h0B51;    16'd29605: out <= 16'h01B1;    16'd29606: out <= 16'hFCF9;    16'd29607: out <= 16'hFEED;
    16'd29608: out <= 16'h090B;    16'd29609: out <= 16'hFB72;    16'd29610: out <= 16'h0772;    16'd29611: out <= 16'h04DE;
    16'd29612: out <= 16'hFF22;    16'd29613: out <= 16'h01CB;    16'd29614: out <= 16'h01DF;    16'd29615: out <= 16'h051E;
    16'd29616: out <= 16'h018C;    16'd29617: out <= 16'h0022;    16'd29618: out <= 16'h0656;    16'd29619: out <= 16'h05AD;
    16'd29620: out <= 16'h094E;    16'd29621: out <= 16'h0B54;    16'd29622: out <= 16'hFF94;    16'd29623: out <= 16'h0B75;
    16'd29624: out <= 16'h0927;    16'd29625: out <= 16'hFC3A;    16'd29626: out <= 16'h04D5;    16'd29627: out <= 16'hFFA7;
    16'd29628: out <= 16'hFE16;    16'd29629: out <= 16'h01DE;    16'd29630: out <= 16'h05F9;    16'd29631: out <= 16'h05EF;
    16'd29632: out <= 16'h0318;    16'd29633: out <= 16'h0559;    16'd29634: out <= 16'h02CA;    16'd29635: out <= 16'h02A5;
    16'd29636: out <= 16'h01EC;    16'd29637: out <= 16'h07EC;    16'd29638: out <= 16'h02BA;    16'd29639: out <= 16'h0C13;
    16'd29640: out <= 16'h022D;    16'd29641: out <= 16'hFCA4;    16'd29642: out <= 16'h0744;    16'd29643: out <= 16'h0028;
    16'd29644: out <= 16'h0420;    16'd29645: out <= 16'h0764;    16'd29646: out <= 16'h060C;    16'd29647: out <= 16'hFF53;
    16'd29648: out <= 16'h07BE;    16'd29649: out <= 16'h07A2;    16'd29650: out <= 16'hFFD1;    16'd29651: out <= 16'hFE66;
    16'd29652: out <= 16'h03D1;    16'd29653: out <= 16'h03B8;    16'd29654: out <= 16'h0520;    16'd29655: out <= 16'h014E;
    16'd29656: out <= 16'hFC3C;    16'd29657: out <= 16'h0087;    16'd29658: out <= 16'hF930;    16'd29659: out <= 16'hFDF6;
    16'd29660: out <= 16'h042A;    16'd29661: out <= 16'h00B5;    16'd29662: out <= 16'hFEB0;    16'd29663: out <= 16'h0077;
    16'd29664: out <= 16'hFF5E;    16'd29665: out <= 16'h04E0;    16'd29666: out <= 16'h005A;    16'd29667: out <= 16'h0262;
    16'd29668: out <= 16'h010D;    16'd29669: out <= 16'h0152;    16'd29670: out <= 16'h02E2;    16'd29671: out <= 16'h00B0;
    16'd29672: out <= 16'h041E;    16'd29673: out <= 16'hFB10;    16'd29674: out <= 16'h0110;    16'd29675: out <= 16'h0152;
    16'd29676: out <= 16'h0328;    16'd29677: out <= 16'hFAE9;    16'd29678: out <= 16'hF868;    16'd29679: out <= 16'h0090;
    16'd29680: out <= 16'hFCAB;    16'd29681: out <= 16'h0163;    16'd29682: out <= 16'h03C7;    16'd29683: out <= 16'hFF28;
    16'd29684: out <= 16'h087D;    16'd29685: out <= 16'hFC07;    16'd29686: out <= 16'hFAAD;    16'd29687: out <= 16'h0177;
    16'd29688: out <= 16'h0392;    16'd29689: out <= 16'hFAA3;    16'd29690: out <= 16'h023F;    16'd29691: out <= 16'h07A9;
    16'd29692: out <= 16'h00DE;    16'd29693: out <= 16'h0492;    16'd29694: out <= 16'hFF50;    16'd29695: out <= 16'hFDF3;
    16'd29696: out <= 16'h02CB;    16'd29697: out <= 16'h02F6;    16'd29698: out <= 16'h012F;    16'd29699: out <= 16'hFB1D;
    16'd29700: out <= 16'hFF93;    16'd29701: out <= 16'hFD1A;    16'd29702: out <= 16'h0018;    16'd29703: out <= 16'hFB2F;
    16'd29704: out <= 16'hFD7B;    16'd29705: out <= 16'h01D7;    16'd29706: out <= 16'hFCE5;    16'd29707: out <= 16'h0610;
    16'd29708: out <= 16'h0179;    16'd29709: out <= 16'h007E;    16'd29710: out <= 16'hFBE3;    16'd29711: out <= 16'hFB6E;
    16'd29712: out <= 16'hFD53;    16'd29713: out <= 16'hF960;    16'd29714: out <= 16'h0281;    16'd29715: out <= 16'hFCE0;
    16'd29716: out <= 16'h048D;    16'd29717: out <= 16'hFB92;    16'd29718: out <= 16'hFB67;    16'd29719: out <= 16'h0355;
    16'd29720: out <= 16'h0B5F;    16'd29721: out <= 16'hFE4D;    16'd29722: out <= 16'h057E;    16'd29723: out <= 16'h03A3;
    16'd29724: out <= 16'h02C2;    16'd29725: out <= 16'h0775;    16'd29726: out <= 16'h06DF;    16'd29727: out <= 16'h0373;
    16'd29728: out <= 16'h036B;    16'd29729: out <= 16'h01DF;    16'd29730: out <= 16'h0871;    16'd29731: out <= 16'h0480;
    16'd29732: out <= 16'h0452;    16'd29733: out <= 16'hFFE8;    16'd29734: out <= 16'h0912;    16'd29735: out <= 16'h02FF;
    16'd29736: out <= 16'h0584;    16'd29737: out <= 16'hFE25;    16'd29738: out <= 16'h0525;    16'd29739: out <= 16'h0977;
    16'd29740: out <= 16'hFA75;    16'd29741: out <= 16'h00B5;    16'd29742: out <= 16'h095B;    16'd29743: out <= 16'h02ED;
    16'd29744: out <= 16'h03E9;    16'd29745: out <= 16'h071B;    16'd29746: out <= 16'h0AA5;    16'd29747: out <= 16'h0C9D;
    16'd29748: out <= 16'h0691;    16'd29749: out <= 16'h0724;    16'd29750: out <= 16'h031E;    16'd29751: out <= 16'h038B;
    16'd29752: out <= 16'h0BB1;    16'd29753: out <= 16'h08A9;    16'd29754: out <= 16'h0064;    16'd29755: out <= 16'h0948;
    16'd29756: out <= 16'h0614;    16'd29757: out <= 16'hFF42;    16'd29758: out <= 16'h09E1;    16'd29759: out <= 16'h0849;
    16'd29760: out <= 16'h03C6;    16'd29761: out <= 16'h054A;    16'd29762: out <= 16'hFE95;    16'd29763: out <= 16'hFF10;
    16'd29764: out <= 16'h08D5;    16'd29765: out <= 16'h089C;    16'd29766: out <= 16'h0271;    16'd29767: out <= 16'h0754;
    16'd29768: out <= 16'h0019;    16'd29769: out <= 16'h00E3;    16'd29770: out <= 16'h017D;    16'd29771: out <= 16'hFF5F;
    16'd29772: out <= 16'h01FE;    16'd29773: out <= 16'h00FE;    16'd29774: out <= 16'h0151;    16'd29775: out <= 16'hFEED;
    16'd29776: out <= 16'h0088;    16'd29777: out <= 16'h02B9;    16'd29778: out <= 16'h04C3;    16'd29779: out <= 16'h0226;
    16'd29780: out <= 16'hFC5E;    16'd29781: out <= 16'h09F1;    16'd29782: out <= 16'h018E;    16'd29783: out <= 16'h0C30;
    16'd29784: out <= 16'h0B6B;    16'd29785: out <= 16'hFF25;    16'd29786: out <= 16'h00BB;    16'd29787: out <= 16'h01B2;
    16'd29788: out <= 16'hFD67;    16'd29789: out <= 16'hF9E0;    16'd29790: out <= 16'h0241;    16'd29791: out <= 16'h0516;
    16'd29792: out <= 16'h00CB;    16'd29793: out <= 16'h04A2;    16'd29794: out <= 16'h039B;    16'd29795: out <= 16'h0C57;
    16'd29796: out <= 16'h0573;    16'd29797: out <= 16'hFEB5;    16'd29798: out <= 16'h00F1;    16'd29799: out <= 16'h0684;
    16'd29800: out <= 16'h03A4;    16'd29801: out <= 16'h0195;    16'd29802: out <= 16'h0003;    16'd29803: out <= 16'hFD85;
    16'd29804: out <= 16'hFF2B;    16'd29805: out <= 16'hF9CA;    16'd29806: out <= 16'hFEDA;    16'd29807: out <= 16'h0B2B;
    16'd29808: out <= 16'h0058;    16'd29809: out <= 16'hFDCE;    16'd29810: out <= 16'h0211;    16'd29811: out <= 16'h02B1;
    16'd29812: out <= 16'h03CA;    16'd29813: out <= 16'h040E;    16'd29814: out <= 16'hFF5A;    16'd29815: out <= 16'h0367;
    16'd29816: out <= 16'h01BC;    16'd29817: out <= 16'h0521;    16'd29818: out <= 16'hFCED;    16'd29819: out <= 16'h0030;
    16'd29820: out <= 16'h0482;    16'd29821: out <= 16'h04DF;    16'd29822: out <= 16'h045A;    16'd29823: out <= 16'h0331;
    16'd29824: out <= 16'h0B3A;    16'd29825: out <= 16'hFD4F;    16'd29826: out <= 16'h072E;    16'd29827: out <= 16'h05D0;
    16'd29828: out <= 16'h0226;    16'd29829: out <= 16'h0313;    16'd29830: out <= 16'h062C;    16'd29831: out <= 16'h0066;
    16'd29832: out <= 16'h0587;    16'd29833: out <= 16'h07BB;    16'd29834: out <= 16'h005C;    16'd29835: out <= 16'h0129;
    16'd29836: out <= 16'h02FA;    16'd29837: out <= 16'h0998;    16'd29838: out <= 16'h0571;    16'd29839: out <= 16'h014C;
    16'd29840: out <= 16'h06BC;    16'd29841: out <= 16'h03AF;    16'd29842: out <= 16'h00BE;    16'd29843: out <= 16'hFF23;
    16'd29844: out <= 16'h0398;    16'd29845: out <= 16'h0374;    16'd29846: out <= 16'h07EA;    16'd29847: out <= 16'hFF15;
    16'd29848: out <= 16'h04D7;    16'd29849: out <= 16'h0846;    16'd29850: out <= 16'h08CA;    16'd29851: out <= 16'h068A;
    16'd29852: out <= 16'h05E4;    16'd29853: out <= 16'h0C5C;    16'd29854: out <= 16'hFF50;    16'd29855: out <= 16'h0742;
    16'd29856: out <= 16'h05F0;    16'd29857: out <= 16'h0362;    16'd29858: out <= 16'h0259;    16'd29859: out <= 16'hFC66;
    16'd29860: out <= 16'h02BC;    16'd29861: out <= 16'h0630;    16'd29862: out <= 16'hFD84;    16'd29863: out <= 16'h054C;
    16'd29864: out <= 16'hFE76;    16'd29865: out <= 16'h01CF;    16'd29866: out <= 16'hFE09;    16'd29867: out <= 16'h03AA;
    16'd29868: out <= 16'h0426;    16'd29869: out <= 16'h0374;    16'd29870: out <= 16'hFF9A;    16'd29871: out <= 16'h06EE;
    16'd29872: out <= 16'h073F;    16'd29873: out <= 16'hFF50;    16'd29874: out <= 16'h0079;    16'd29875: out <= 16'h05EB;
    16'd29876: out <= 16'h08E7;    16'd29877: out <= 16'h056B;    16'd29878: out <= 16'h0219;    16'd29879: out <= 16'h0518;
    16'd29880: out <= 16'hFEC1;    16'd29881: out <= 16'h028E;    16'd29882: out <= 16'h05DC;    16'd29883: out <= 16'h00D2;
    16'd29884: out <= 16'hFFCF;    16'd29885: out <= 16'h0369;    16'd29886: out <= 16'h022D;    16'd29887: out <= 16'h00AD;
    16'd29888: out <= 16'h0B8A;    16'd29889: out <= 16'h060E;    16'd29890: out <= 16'hFF22;    16'd29891: out <= 16'h0313;
    16'd29892: out <= 16'h0800;    16'd29893: out <= 16'h0701;    16'd29894: out <= 16'h0060;    16'd29895: out <= 16'h055E;
    16'd29896: out <= 16'h05C9;    16'd29897: out <= 16'hFF63;    16'd29898: out <= 16'h06B1;    16'd29899: out <= 16'h054D;
    16'd29900: out <= 16'h0962;    16'd29901: out <= 16'h049F;    16'd29902: out <= 16'h06D1;    16'd29903: out <= 16'h0310;
    16'd29904: out <= 16'h07D5;    16'd29905: out <= 16'h026C;    16'd29906: out <= 16'h02EA;    16'd29907: out <= 16'h03C6;
    16'd29908: out <= 16'h09B5;    16'd29909: out <= 16'hFE99;    16'd29910: out <= 16'h054E;    16'd29911: out <= 16'h0751;
    16'd29912: out <= 16'h0482;    16'd29913: out <= 16'h003D;    16'd29914: out <= 16'hFC37;    16'd29915: out <= 16'h06C2;
    16'd29916: out <= 16'h0505;    16'd29917: out <= 16'h0116;    16'd29918: out <= 16'h0035;    16'd29919: out <= 16'h012A;
    16'd29920: out <= 16'h07A6;    16'd29921: out <= 16'h010F;    16'd29922: out <= 16'h0402;    16'd29923: out <= 16'h01BD;
    16'd29924: out <= 16'h0A88;    16'd29925: out <= 16'hF67D;    16'd29926: out <= 16'h03B4;    16'd29927: out <= 16'h043F;
    16'd29928: out <= 16'h049C;    16'd29929: out <= 16'hFD73;    16'd29930: out <= 16'hFB4B;    16'd29931: out <= 16'h0139;
    16'd29932: out <= 16'hFDFF;    16'd29933: out <= 16'hFF75;    16'd29934: out <= 16'hFEEE;    16'd29935: out <= 16'h01D4;
    16'd29936: out <= 16'hF747;    16'd29937: out <= 16'h01C9;    16'd29938: out <= 16'hFC3C;    16'd29939: out <= 16'hFDD0;
    16'd29940: out <= 16'h01F4;    16'd29941: out <= 16'h008E;    16'd29942: out <= 16'hFF51;    16'd29943: out <= 16'hFF1A;
    16'd29944: out <= 16'hFD70;    16'd29945: out <= 16'h06C5;    16'd29946: out <= 16'h04FF;    16'd29947: out <= 16'h010D;
    16'd29948: out <= 16'hFD69;    16'd29949: out <= 16'h00B6;    16'd29950: out <= 16'h0102;    16'd29951: out <= 16'h087A;
    16'd29952: out <= 16'h03B3;    16'd29953: out <= 16'h0398;    16'd29954: out <= 16'h016C;    16'd29955: out <= 16'h043F;
    16'd29956: out <= 16'hFB88;    16'd29957: out <= 16'h01AB;    16'd29958: out <= 16'h01E3;    16'd29959: out <= 16'h0561;
    16'd29960: out <= 16'h0341;    16'd29961: out <= 16'hF826;    16'd29962: out <= 16'hFE54;    16'd29963: out <= 16'h01D9;
    16'd29964: out <= 16'hFA79;    16'd29965: out <= 16'hFF4E;    16'd29966: out <= 16'hFB8E;    16'd29967: out <= 16'h0531;
    16'd29968: out <= 16'h052D;    16'd29969: out <= 16'h030A;    16'd29970: out <= 16'h07D5;    16'd29971: out <= 16'hFF9E;
    16'd29972: out <= 16'h0434;    16'd29973: out <= 16'hF7A7;    16'd29974: out <= 16'h05C6;    16'd29975: out <= 16'h09C1;
    16'd29976: out <= 16'h04A0;    16'd29977: out <= 16'hF7E8;    16'd29978: out <= 16'h0372;    16'd29979: out <= 16'h040D;
    16'd29980: out <= 16'h026B;    16'd29981: out <= 16'h05AD;    16'd29982: out <= 16'h0409;    16'd29983: out <= 16'h0297;
    16'd29984: out <= 16'h03ED;    16'd29985: out <= 16'hFD7C;    16'd29986: out <= 16'h08BF;    16'd29987: out <= 16'hFEF2;
    16'd29988: out <= 16'hFFE2;    16'd29989: out <= 16'h0441;    16'd29990: out <= 16'h0077;    16'd29991: out <= 16'h0764;
    16'd29992: out <= 16'h05CA;    16'd29993: out <= 16'h022E;    16'd29994: out <= 16'h016C;    16'd29995: out <= 16'h060D;
    16'd29996: out <= 16'h01AF;    16'd29997: out <= 16'h06FA;    16'd29998: out <= 16'h07D0;    16'd29999: out <= 16'hFF2C;
    16'd30000: out <= 16'h07D3;    16'd30001: out <= 16'hFB58;    16'd30002: out <= 16'h02E5;    16'd30003: out <= 16'h03FE;
    16'd30004: out <= 16'h090F;    16'd30005: out <= 16'h044A;    16'd30006: out <= 16'h0906;    16'd30007: out <= 16'hFC2F;
    16'd30008: out <= 16'hFB44;    16'd30009: out <= 16'h0617;    16'd30010: out <= 16'h0597;    16'd30011: out <= 16'h04A1;
    16'd30012: out <= 16'h0B8B;    16'd30013: out <= 16'h04C8;    16'd30014: out <= 16'h091D;    16'd30015: out <= 16'h014A;
    16'd30016: out <= 16'h03BA;    16'd30017: out <= 16'h0060;    16'd30018: out <= 16'h0737;    16'd30019: out <= 16'hFBF9;
    16'd30020: out <= 16'h0114;    16'd30021: out <= 16'h0702;    16'd30022: out <= 16'h0774;    16'd30023: out <= 16'h05CE;
    16'd30024: out <= 16'h026F;    16'd30025: out <= 16'h0940;    16'd30026: out <= 16'h0148;    16'd30027: out <= 16'h04DC;
    16'd30028: out <= 16'h0858;    16'd30029: out <= 16'hFDE8;    16'd30030: out <= 16'h066D;    16'd30031: out <= 16'h004F;
    16'd30032: out <= 16'hFFA9;    16'd30033: out <= 16'h04A1;    16'd30034: out <= 16'h060E;    16'd30035: out <= 16'h04B7;
    16'd30036: out <= 16'h05C5;    16'd30037: out <= 16'hFFF8;    16'd30038: out <= 16'h058E;    16'd30039: out <= 16'h0324;
    16'd30040: out <= 16'h055C;    16'd30041: out <= 16'h098A;    16'd30042: out <= 16'h05AA;    16'd30043: out <= 16'h043C;
    16'd30044: out <= 16'h07AF;    16'd30045: out <= 16'h01F8;    16'd30046: out <= 16'h0428;    16'd30047: out <= 16'h080B;
    16'd30048: out <= 16'h098B;    16'd30049: out <= 16'h0375;    16'd30050: out <= 16'hFFFC;    16'd30051: out <= 16'h0796;
    16'd30052: out <= 16'h0273;    16'd30053: out <= 16'h05F6;    16'd30054: out <= 16'h0411;    16'd30055: out <= 16'h01BF;
    16'd30056: out <= 16'hFD52;    16'd30057: out <= 16'hFD79;    16'd30058: out <= 16'h02BF;    16'd30059: out <= 16'h06DF;
    16'd30060: out <= 16'h06C0;    16'd30061: out <= 16'h0A05;    16'd30062: out <= 16'h07A7;    16'd30063: out <= 16'h06D8;
    16'd30064: out <= 16'h01A8;    16'd30065: out <= 16'h0717;    16'd30066: out <= 16'h01A2;    16'd30067: out <= 16'hFE71;
    16'd30068: out <= 16'h0484;    16'd30069: out <= 16'h0935;    16'd30070: out <= 16'hFFE6;    16'd30071: out <= 16'h0206;
    16'd30072: out <= 16'h0599;    16'd30073: out <= 16'h06B3;    16'd30074: out <= 16'hFE39;    16'd30075: out <= 16'h0458;
    16'd30076: out <= 16'h050B;    16'd30077: out <= 16'h05CB;    16'd30078: out <= 16'hFF97;    16'd30079: out <= 16'h03E4;
    16'd30080: out <= 16'h0099;    16'd30081: out <= 16'h0485;    16'd30082: out <= 16'h009F;    16'd30083: out <= 16'h03C7;
    16'd30084: out <= 16'h044B;    16'd30085: out <= 16'h09D9;    16'd30086: out <= 16'hFFF2;    16'd30087: out <= 16'h0A5C;
    16'd30088: out <= 16'h07A8;    16'd30089: out <= 16'h042E;    16'd30090: out <= 16'h0643;    16'd30091: out <= 16'hFEDA;
    16'd30092: out <= 16'h05DA;    16'd30093: out <= 16'h00B7;    16'd30094: out <= 16'h0166;    16'd30095: out <= 16'h02E0;
    16'd30096: out <= 16'hFE51;    16'd30097: out <= 16'h014F;    16'd30098: out <= 16'h0061;    16'd30099: out <= 16'h0B36;
    16'd30100: out <= 16'h02AB;    16'd30101: out <= 16'h0419;    16'd30102: out <= 16'h032F;    16'd30103: out <= 16'h074A;
    16'd30104: out <= 16'h03B9;    16'd30105: out <= 16'h09F1;    16'd30106: out <= 16'h0683;    16'd30107: out <= 16'h06E0;
    16'd30108: out <= 16'h023C;    16'd30109: out <= 16'h020B;    16'd30110: out <= 16'h0100;    16'd30111: out <= 16'h0384;
    16'd30112: out <= 16'h00E1;    16'd30113: out <= 16'h0567;    16'd30114: out <= 16'h0727;    16'd30115: out <= 16'h05AC;
    16'd30116: out <= 16'h02BB;    16'd30117: out <= 16'h079D;    16'd30118: out <= 16'h0414;    16'd30119: out <= 16'h0168;
    16'd30120: out <= 16'h037C;    16'd30121: out <= 16'h0658;    16'd30122: out <= 16'h0248;    16'd30123: out <= 16'h04D0;
    16'd30124: out <= 16'h00FB;    16'd30125: out <= 16'h0230;    16'd30126: out <= 16'h037E;    16'd30127: out <= 16'h0A15;
    16'd30128: out <= 16'hFD9D;    16'd30129: out <= 16'h07BF;    16'd30130: out <= 16'h010D;    16'd30131: out <= 16'h02AF;
    16'd30132: out <= 16'h04B1;    16'd30133: out <= 16'h092A;    16'd30134: out <= 16'h01D2;    16'd30135: out <= 16'h05C2;
    16'd30136: out <= 16'h0370;    16'd30137: out <= 16'h06E1;    16'd30138: out <= 16'h034D;    16'd30139: out <= 16'h0D55;
    16'd30140: out <= 16'h043D;    16'd30141: out <= 16'h0180;    16'd30142: out <= 16'hFEC2;    16'd30143: out <= 16'h03A0;
    16'd30144: out <= 16'hFD59;    16'd30145: out <= 16'h0048;    16'd30146: out <= 16'h015C;    16'd30147: out <= 16'h0659;
    16'd30148: out <= 16'h009A;    16'd30149: out <= 16'h06C1;    16'd30150: out <= 16'hFD7A;    16'd30151: out <= 16'hFFF7;
    16'd30152: out <= 16'h09FA;    16'd30153: out <= 16'hFBB9;    16'd30154: out <= 16'h076E;    16'd30155: out <= 16'h059C;
    16'd30156: out <= 16'h0189;    16'd30157: out <= 16'h0082;    16'd30158: out <= 16'hFCE9;    16'd30159: out <= 16'hFD6D;
    16'd30160: out <= 16'h0986;    16'd30161: out <= 16'h046B;    16'd30162: out <= 16'hFCC8;    16'd30163: out <= 16'h01C1;
    16'd30164: out <= 16'h0659;    16'd30165: out <= 16'h0677;    16'd30166: out <= 16'h031F;    16'd30167: out <= 16'hFCC4;
    16'd30168: out <= 16'h00AF;    16'd30169: out <= 16'h02B7;    16'd30170: out <= 16'h0708;    16'd30171: out <= 16'hFA69;
    16'd30172: out <= 16'h0459;    16'd30173: out <= 16'h003B;    16'd30174: out <= 16'hFA29;    16'd30175: out <= 16'hF2FA;
    16'd30176: out <= 16'h05C8;    16'd30177: out <= 16'hFECD;    16'd30178: out <= 16'h014F;    16'd30179: out <= 16'h015B;
    16'd30180: out <= 16'h010A;    16'd30181: out <= 16'h00B0;    16'd30182: out <= 16'hFD3C;    16'd30183: out <= 16'hFE00;
    16'd30184: out <= 16'h02BA;    16'd30185: out <= 16'h03AA;    16'd30186: out <= 16'h01CF;    16'd30187: out <= 16'hFBB7;
    16'd30188: out <= 16'h080F;    16'd30189: out <= 16'hF5F7;    16'd30190: out <= 16'hFBE2;    16'd30191: out <= 16'h0208;
    16'd30192: out <= 16'h019A;    16'd30193: out <= 16'h01B3;    16'd30194: out <= 16'hFD62;    16'd30195: out <= 16'hFFA8;
    16'd30196: out <= 16'hFBB9;    16'd30197: out <= 16'hFCF7;    16'd30198: out <= 16'h021B;    16'd30199: out <= 16'hFB82;
    16'd30200: out <= 16'hFCE6;    16'd30201: out <= 16'h05C4;    16'd30202: out <= 16'hFF8F;    16'd30203: out <= 16'h0459;
    16'd30204: out <= 16'h0003;    16'd30205: out <= 16'h06DF;    16'd30206: out <= 16'hFEF8;    16'd30207: out <= 16'h00FD;
    16'd30208: out <= 16'h011E;    16'd30209: out <= 16'hFF08;    16'd30210: out <= 16'h0260;    16'd30211: out <= 16'h0252;
    16'd30212: out <= 16'h06A0;    16'd30213: out <= 16'hFC51;    16'd30214: out <= 16'h0055;    16'd30215: out <= 16'hFCF2;
    16'd30216: out <= 16'h035D;    16'd30217: out <= 16'hFCFC;    16'd30218: out <= 16'hFD8C;    16'd30219: out <= 16'hFEA0;
    16'd30220: out <= 16'h028A;    16'd30221: out <= 16'hFEE2;    16'd30222: out <= 16'h044D;    16'd30223: out <= 16'hFF53;
    16'd30224: out <= 16'h041E;    16'd30225: out <= 16'hF8AF;    16'd30226: out <= 16'hFF01;    16'd30227: out <= 16'hF59F;
    16'd30228: out <= 16'h0187;    16'd30229: out <= 16'hFF90;    16'd30230: out <= 16'h04A1;    16'd30231: out <= 16'h09D6;
    16'd30232: out <= 16'h0037;    16'd30233: out <= 16'h0076;    16'd30234: out <= 16'h036D;    16'd30235: out <= 16'h0ACC;
    16'd30236: out <= 16'h0171;    16'd30237: out <= 16'h03CC;    16'd30238: out <= 16'h0668;    16'd30239: out <= 16'h03D4;
    16'd30240: out <= 16'h06B0;    16'd30241: out <= 16'h095A;    16'd30242: out <= 16'h09FF;    16'd30243: out <= 16'h0287;
    16'd30244: out <= 16'h0612;    16'd30245: out <= 16'h097C;    16'd30246: out <= 16'hFDE9;    16'd30247: out <= 16'h03E7;
    16'd30248: out <= 16'h05DA;    16'd30249: out <= 16'hF9E0;    16'd30250: out <= 16'h096F;    16'd30251: out <= 16'hF860;
    16'd30252: out <= 16'h00A0;    16'd30253: out <= 16'hFF1D;    16'd30254: out <= 16'h0577;    16'd30255: out <= 16'h0782;
    16'd30256: out <= 16'h07E7;    16'd30257: out <= 16'h019E;    16'd30258: out <= 16'h09BB;    16'd30259: out <= 16'h0678;
    16'd30260: out <= 16'h0457;    16'd30261: out <= 16'h0428;    16'd30262: out <= 16'h079A;    16'd30263: out <= 16'h0A66;
    16'd30264: out <= 16'h0758;    16'd30265: out <= 16'h0895;    16'd30266: out <= 16'h07B4;    16'd30267: out <= 16'hFDE7;
    16'd30268: out <= 16'hFFCA;    16'd30269: out <= 16'h00B0;    16'd30270: out <= 16'h0931;    16'd30271: out <= 16'h02D8;
    16'd30272: out <= 16'h0625;    16'd30273: out <= 16'h06E4;    16'd30274: out <= 16'h04B8;    16'd30275: out <= 16'hFDE4;
    16'd30276: out <= 16'h0268;    16'd30277: out <= 16'h0283;    16'd30278: out <= 16'h07D0;    16'd30279: out <= 16'h0634;
    16'd30280: out <= 16'h0654;    16'd30281: out <= 16'hFE1E;    16'd30282: out <= 16'h04FD;    16'd30283: out <= 16'h05D0;
    16'd30284: out <= 16'h02AC;    16'd30285: out <= 16'h0921;    16'd30286: out <= 16'h02B4;    16'd30287: out <= 16'hFBD3;
    16'd30288: out <= 16'h011C;    16'd30289: out <= 16'h04CA;    16'd30290: out <= 16'hFED3;    16'd30291: out <= 16'h0247;
    16'd30292: out <= 16'h05DE;    16'd30293: out <= 16'h03FB;    16'd30294: out <= 16'h0AD4;    16'd30295: out <= 16'h0332;
    16'd30296: out <= 16'h02FD;    16'd30297: out <= 16'h01FE;    16'd30298: out <= 16'h0363;    16'd30299: out <= 16'h076D;
    16'd30300: out <= 16'h0225;    16'd30301: out <= 16'h02D9;    16'd30302: out <= 16'h0320;    16'd30303: out <= 16'hFFD0;
    16'd30304: out <= 16'h0378;    16'd30305: out <= 16'h0E58;    16'd30306: out <= 16'h048F;    16'd30307: out <= 16'hFD73;
    16'd30308: out <= 16'h01C2;    16'd30309: out <= 16'h0390;    16'd30310: out <= 16'h01B6;    16'd30311: out <= 16'h0299;
    16'd30312: out <= 16'h0988;    16'd30313: out <= 16'h06DF;    16'd30314: out <= 16'h025C;    16'd30315: out <= 16'h0B5D;
    16'd30316: out <= 16'h0619;    16'd30317: out <= 16'h0555;    16'd30318: out <= 16'h0683;    16'd30319: out <= 16'hFFA2;
    16'd30320: out <= 16'h06B1;    16'd30321: out <= 16'h049C;    16'd30322: out <= 16'h028C;    16'd30323: out <= 16'h032B;
    16'd30324: out <= 16'h0743;    16'd30325: out <= 16'h04FA;    16'd30326: out <= 16'h06AD;    16'd30327: out <= 16'h020E;
    16'd30328: out <= 16'h0279;    16'd30329: out <= 16'h0030;    16'd30330: out <= 16'h00D4;    16'd30331: out <= 16'h02AF;
    16'd30332: out <= 16'h07A8;    16'd30333: out <= 16'h008A;    16'd30334: out <= 16'h0002;    16'd30335: out <= 16'h0498;
    16'd30336: out <= 16'hFF82;    16'd30337: out <= 16'h0149;    16'd30338: out <= 16'h06E6;    16'd30339: out <= 16'h00BC;
    16'd30340: out <= 16'hFFB8;    16'd30341: out <= 16'h08C3;    16'd30342: out <= 16'h0633;    16'd30343: out <= 16'h08B4;
    16'd30344: out <= 16'h04ED;    16'd30345: out <= 16'h041A;    16'd30346: out <= 16'h02EC;    16'd30347: out <= 16'h03AE;
    16'd30348: out <= 16'h084F;    16'd30349: out <= 16'h05E3;    16'd30350: out <= 16'h0458;    16'd30351: out <= 16'h09CE;
    16'd30352: out <= 16'h06C4;    16'd30353: out <= 16'h08F1;    16'd30354: out <= 16'h075C;    16'd30355: out <= 16'h01F3;
    16'd30356: out <= 16'hFE50;    16'd30357: out <= 16'h00EA;    16'd30358: out <= 16'h0BD0;    16'd30359: out <= 16'h05AC;
    16'd30360: out <= 16'h084D;    16'd30361: out <= 16'h0278;    16'd30362: out <= 16'h04AD;    16'd30363: out <= 16'h04C0;
    16'd30364: out <= 16'hFF37;    16'd30365: out <= 16'h0909;    16'd30366: out <= 16'h02B5;    16'd30367: out <= 16'h0183;
    16'd30368: out <= 16'hFDCF;    16'd30369: out <= 16'h0733;    16'd30370: out <= 16'h0564;    16'd30371: out <= 16'h0292;
    16'd30372: out <= 16'h0971;    16'd30373: out <= 16'h011F;    16'd30374: out <= 16'hFE50;    16'd30375: out <= 16'h05C4;
    16'd30376: out <= 16'hFD00;    16'd30377: out <= 16'h0557;    16'd30378: out <= 16'h0BD2;    16'd30379: out <= 16'h03B0;
    16'd30380: out <= 16'h0073;    16'd30381: out <= 16'h05A7;    16'd30382: out <= 16'hFDB3;    16'd30383: out <= 16'h0460;
    16'd30384: out <= 16'h0573;    16'd30385: out <= 16'h0C51;    16'd30386: out <= 16'h0A0D;    16'd30387: out <= 16'h0A28;
    16'd30388: out <= 16'h09A5;    16'd30389: out <= 16'h0723;    16'd30390: out <= 16'h0569;    16'd30391: out <= 16'h0385;
    16'd30392: out <= 16'h0723;    16'd30393: out <= 16'hFFC7;    16'd30394: out <= 16'hFEB4;    16'd30395: out <= 16'hFC47;
    16'd30396: out <= 16'hFFFB;    16'd30397: out <= 16'h0E88;    16'd30398: out <= 16'h0891;    16'd30399: out <= 16'h05A5;
    16'd30400: out <= 16'h0576;    16'd30401: out <= 16'h062A;    16'd30402: out <= 16'h05CF;    16'd30403: out <= 16'hFEED;
    16'd30404: out <= 16'h05B8;    16'd30405: out <= 16'h0254;    16'd30406: out <= 16'h06CA;    16'd30407: out <= 16'h0380;
    16'd30408: out <= 16'h0110;    16'd30409: out <= 16'h03F6;    16'd30410: out <= 16'h0397;    16'd30411: out <= 16'h038A;
    16'd30412: out <= 16'h0791;    16'd30413: out <= 16'h033F;    16'd30414: out <= 16'h06BF;    16'd30415: out <= 16'hFEDD;
    16'd30416: out <= 16'h0491;    16'd30417: out <= 16'hFCCE;    16'd30418: out <= 16'hFFBD;    16'd30419: out <= 16'h0385;
    16'd30420: out <= 16'h0B9B;    16'd30421: out <= 16'hFB70;    16'd30422: out <= 16'h037B;    16'd30423: out <= 16'h05FB;
    16'd30424: out <= 16'hFEC8;    16'd30425: out <= 16'h04B4;    16'd30426: out <= 16'hFC56;    16'd30427: out <= 16'hFD47;
    16'd30428: out <= 16'h009D;    16'd30429: out <= 16'h045E;    16'd30430: out <= 16'hFF25;    16'd30431: out <= 16'hFB5D;
    16'd30432: out <= 16'h02DD;    16'd30433: out <= 16'h0178;    16'd30434: out <= 16'hFD06;    16'd30435: out <= 16'h0190;
    16'd30436: out <= 16'h024B;    16'd30437: out <= 16'h07CD;    16'd30438: out <= 16'hFBE4;    16'd30439: out <= 16'h0250;
    16'd30440: out <= 16'h0855;    16'd30441: out <= 16'hFF73;    16'd30442: out <= 16'hFE60;    16'd30443: out <= 16'hFF96;
    16'd30444: out <= 16'hFCE1;    16'd30445: out <= 16'hFC25;    16'd30446: out <= 16'hFA1B;    16'd30447: out <= 16'h05D4;
    16'd30448: out <= 16'h00E7;    16'd30449: out <= 16'hFF8D;    16'd30450: out <= 16'h097A;    16'd30451: out <= 16'hFDAA;
    16'd30452: out <= 16'h0493;    16'd30453: out <= 16'hFDA9;    16'd30454: out <= 16'h00D1;    16'd30455: out <= 16'hFB73;
    16'd30456: out <= 16'hFC90;    16'd30457: out <= 16'h03C9;    16'd30458: out <= 16'hFE71;    16'd30459: out <= 16'hFF7A;
    16'd30460: out <= 16'hFBD9;    16'd30461: out <= 16'hFC85;    16'd30462: out <= 16'hFDC5;    16'd30463: out <= 16'hFBBD;
    16'd30464: out <= 16'hFD2C;    16'd30465: out <= 16'h01A4;    16'd30466: out <= 16'hFC34;    16'd30467: out <= 16'hFE70;
    16'd30468: out <= 16'hFBC3;    16'd30469: out <= 16'hFBED;    16'd30470: out <= 16'hFE08;    16'd30471: out <= 16'hF98D;
    16'd30472: out <= 16'hFD61;    16'd30473: out <= 16'hFB35;    16'd30474: out <= 16'hFE65;    16'd30475: out <= 16'h0560;
    16'd30476: out <= 16'h004F;    16'd30477: out <= 16'hFC6A;    16'd30478: out <= 16'hFAB0;    16'd30479: out <= 16'hF68E;
    16'd30480: out <= 16'hFCE8;    16'd30481: out <= 16'h083C;    16'd30482: out <= 16'h0233;    16'd30483: out <= 16'h00EB;
    16'd30484: out <= 16'h01C1;    16'd30485: out <= 16'h005A;    16'd30486: out <= 16'h0386;    16'd30487: out <= 16'h04B3;
    16'd30488: out <= 16'h07C2;    16'd30489: out <= 16'h094A;    16'd30490: out <= 16'h02D8;    16'd30491: out <= 16'h07B8;
    16'd30492: out <= 16'h0611;    16'd30493: out <= 16'h06F4;    16'd30494: out <= 16'h00B1;    16'd30495: out <= 16'h021F;
    16'd30496: out <= 16'h0434;    16'd30497: out <= 16'hFFA3;    16'd30498: out <= 16'h082B;    16'd30499: out <= 16'hFD6B;
    16'd30500: out <= 16'h06F2;    16'd30501: out <= 16'h02C9;    16'd30502: out <= 16'h0551;    16'd30503: out <= 16'h0178;
    16'd30504: out <= 16'h01F2;    16'd30505: out <= 16'h0628;    16'd30506: out <= 16'h0818;    16'd30507: out <= 16'h0273;
    16'd30508: out <= 16'h023C;    16'd30509: out <= 16'h0C2B;    16'd30510: out <= 16'h049E;    16'd30511: out <= 16'h03F7;
    16'd30512: out <= 16'h0607;    16'd30513: out <= 16'h00FD;    16'd30514: out <= 16'h065B;    16'd30515: out <= 16'h038A;
    16'd30516: out <= 16'h05F8;    16'd30517: out <= 16'h0435;    16'd30518: out <= 16'h05D4;    16'd30519: out <= 16'h071F;
    16'd30520: out <= 16'h06EA;    16'd30521: out <= 16'hFB9F;    16'd30522: out <= 16'h0B25;    16'd30523: out <= 16'h04F9;
    16'd30524: out <= 16'h045D;    16'd30525: out <= 16'h02BF;    16'd30526: out <= 16'hF955;    16'd30527: out <= 16'h01A2;
    16'd30528: out <= 16'hFE26;    16'd30529: out <= 16'h0432;    16'd30530: out <= 16'hFA21;    16'd30531: out <= 16'h02B2;
    16'd30532: out <= 16'h0224;    16'd30533: out <= 16'h00A1;    16'd30534: out <= 16'h0017;    16'd30535: out <= 16'hFAFD;
    16'd30536: out <= 16'h0241;    16'd30537: out <= 16'h0646;    16'd30538: out <= 16'h030E;    16'd30539: out <= 16'h0D31;
    16'd30540: out <= 16'h010C;    16'd30541: out <= 16'h05D6;    16'd30542: out <= 16'h09C9;    16'd30543: out <= 16'hFF96;
    16'd30544: out <= 16'h0785;    16'd30545: out <= 16'h039D;    16'd30546: out <= 16'hFBCC;    16'd30547: out <= 16'hFEF5;
    16'd30548: out <= 16'h00C7;    16'd30549: out <= 16'h0010;    16'd30550: out <= 16'h05A7;    16'd30551: out <= 16'h027D;
    16'd30552: out <= 16'h0646;    16'd30553: out <= 16'h0108;    16'd30554: out <= 16'h0520;    16'd30555: out <= 16'h03B0;
    16'd30556: out <= 16'h0C5D;    16'd30557: out <= 16'h0C76;    16'd30558: out <= 16'h087A;    16'd30559: out <= 16'h086C;
    16'd30560: out <= 16'h0016;    16'd30561: out <= 16'h03D3;    16'd30562: out <= 16'h0793;    16'd30563: out <= 16'h0171;
    16'd30564: out <= 16'h039F;    16'd30565: out <= 16'h08C6;    16'd30566: out <= 16'h0D71;    16'd30567: out <= 16'h013C;
    16'd30568: out <= 16'hFFD0;    16'd30569: out <= 16'hFD68;    16'd30570: out <= 16'h064A;    16'd30571: out <= 16'h08EE;
    16'd30572: out <= 16'hFEEA;    16'd30573: out <= 16'h06D1;    16'd30574: out <= 16'h05EC;    16'd30575: out <= 16'h018E;
    16'd30576: out <= 16'h06B8;    16'd30577: out <= 16'h03AE;    16'd30578: out <= 16'hFD83;    16'd30579: out <= 16'h0763;
    16'd30580: out <= 16'h0D5F;    16'd30581: out <= 16'h009A;    16'd30582: out <= 16'h0B9A;    16'd30583: out <= 16'h05D8;
    16'd30584: out <= 16'h078D;    16'd30585: out <= 16'h0F4D;    16'd30586: out <= 16'h053F;    16'd30587: out <= 16'hFFC4;
    16'd30588: out <= 16'h0460;    16'd30589: out <= 16'h05C9;    16'd30590: out <= 16'h0413;    16'd30591: out <= 16'h0139;
    16'd30592: out <= 16'h02F1;    16'd30593: out <= 16'h07D0;    16'd30594: out <= 16'h04EA;    16'd30595: out <= 16'h02BF;
    16'd30596: out <= 16'h0331;    16'd30597: out <= 16'h00AA;    16'd30598: out <= 16'h040C;    16'd30599: out <= 16'h0A91;
    16'd30600: out <= 16'h02E2;    16'd30601: out <= 16'h066E;    16'd30602: out <= 16'hFDCC;    16'd30603: out <= 16'h03CF;
    16'd30604: out <= 16'h05FD;    16'd30605: out <= 16'h0669;    16'd30606: out <= 16'h05CB;    16'd30607: out <= 16'h0535;
    16'd30608: out <= 16'h09B2;    16'd30609: out <= 16'h07FF;    16'd30610: out <= 16'h0118;    16'd30611: out <= 16'h07DF;
    16'd30612: out <= 16'h00C4;    16'd30613: out <= 16'h0111;    16'd30614: out <= 16'h0386;    16'd30615: out <= 16'h0566;
    16'd30616: out <= 16'h049D;    16'd30617: out <= 16'h02E7;    16'd30618: out <= 16'h081D;    16'd30619: out <= 16'h0559;
    16'd30620: out <= 16'h0977;    16'd30621: out <= 16'h03EE;    16'd30622: out <= 16'h01DA;    16'd30623: out <= 16'h0403;
    16'd30624: out <= 16'h05D5;    16'd30625: out <= 16'hFBE3;    16'd30626: out <= 16'h000E;    16'd30627: out <= 16'h0220;
    16'd30628: out <= 16'h00E2;    16'd30629: out <= 16'h08CD;    16'd30630: out <= 16'h01D4;    16'd30631: out <= 16'hFCE0;
    16'd30632: out <= 16'h0400;    16'd30633: out <= 16'h05D8;    16'd30634: out <= 16'h0431;    16'd30635: out <= 16'h07E9;
    16'd30636: out <= 16'h02F1;    16'd30637: out <= 16'h0437;    16'd30638: out <= 16'h05A8;    16'd30639: out <= 16'h0244;
    16'd30640: out <= 16'h00A2;    16'd30641: out <= 16'h0C75;    16'd30642: out <= 16'h050B;    16'd30643: out <= 16'hFD55;
    16'd30644: out <= 16'hFD2D;    16'd30645: out <= 16'h0A04;    16'd30646: out <= 16'h0495;    16'd30647: out <= 16'h0B56;
    16'd30648: out <= 16'h0729;    16'd30649: out <= 16'h0AC3;    16'd30650: out <= 16'h06AC;    16'd30651: out <= 16'h02B8;
    16'd30652: out <= 16'hFCA2;    16'd30653: out <= 16'h0962;    16'd30654: out <= 16'h03F4;    16'd30655: out <= 16'h033A;
    16'd30656: out <= 16'h0B3F;    16'd30657: out <= 16'h07AA;    16'd30658: out <= 16'hFD84;    16'd30659: out <= 16'h057E;
    16'd30660: out <= 16'h04FA;    16'd30661: out <= 16'h0951;    16'd30662: out <= 16'h054B;    16'd30663: out <= 16'h08FD;
    16'd30664: out <= 16'h05BE;    16'd30665: out <= 16'hFF53;    16'd30666: out <= 16'h08B0;    16'd30667: out <= 16'hFD69;
    16'd30668: out <= 16'h0437;    16'd30669: out <= 16'h0410;    16'd30670: out <= 16'h049A;    16'd30671: out <= 16'hFD26;
    16'd30672: out <= 16'h04BD;    16'd30673: out <= 16'h069A;    16'd30674: out <= 16'h0836;    16'd30675: out <= 16'h0060;
    16'd30676: out <= 16'h053B;    16'd30677: out <= 16'h04D5;    16'd30678: out <= 16'h0872;    16'd30679: out <= 16'h0170;
    16'd30680: out <= 16'h0330;    16'd30681: out <= 16'hFFDE;    16'd30682: out <= 16'h033B;    16'd30683: out <= 16'h08F1;
    16'd30684: out <= 16'hFE48;    16'd30685: out <= 16'hFDDE;    16'd30686: out <= 16'h02B9;    16'd30687: out <= 16'hFB83;
    16'd30688: out <= 16'h023D;    16'd30689: out <= 16'h08A0;    16'd30690: out <= 16'hFD4E;    16'd30691: out <= 16'h0112;
    16'd30692: out <= 16'hFE96;    16'd30693: out <= 16'h01BE;    16'd30694: out <= 16'h07C7;    16'd30695: out <= 16'h05D9;
    16'd30696: out <= 16'h0034;    16'd30697: out <= 16'h03BE;    16'd30698: out <= 16'hFE72;    16'd30699: out <= 16'hFBB5;
    16'd30700: out <= 16'hFF9E;    16'd30701: out <= 16'hFFC1;    16'd30702: out <= 16'hFC3E;    16'd30703: out <= 16'h0129;
    16'd30704: out <= 16'hFED4;    16'd30705: out <= 16'hFCE6;    16'd30706: out <= 16'h03A1;    16'd30707: out <= 16'hFE28;
    16'd30708: out <= 16'h0114;    16'd30709: out <= 16'hFAF5;    16'd30710: out <= 16'h01AC;    16'd30711: out <= 16'hFFEC;
    16'd30712: out <= 16'h0196;    16'd30713: out <= 16'h057B;    16'd30714: out <= 16'hFD9F;    16'd30715: out <= 16'h0543;
    16'd30716: out <= 16'h0329;    16'd30717: out <= 16'hF9CC;    16'd30718: out <= 16'hF87A;    16'd30719: out <= 16'h04F3;
    16'd30720: out <= 16'hFE84;    16'd30721: out <= 16'h00D4;    16'd30722: out <= 16'hFBFA;    16'd30723: out <= 16'h06DC;
    16'd30724: out <= 16'h004A;    16'd30725: out <= 16'h0112;    16'd30726: out <= 16'hFC0B;    16'd30727: out <= 16'hFFAA;
    16'd30728: out <= 16'h02BA;    16'd30729: out <= 16'h039A;    16'd30730: out <= 16'hF917;    16'd30731: out <= 16'h02D2;
    16'd30732: out <= 16'h0158;    16'd30733: out <= 16'h030B;    16'd30734: out <= 16'hFA2F;    16'd30735: out <= 16'h0660;
    16'd30736: out <= 16'hFF86;    16'd30737: out <= 16'h014F;    16'd30738: out <= 16'hFDA0;    16'd30739: out <= 16'hFDC1;
    16'd30740: out <= 16'h0150;    16'd30741: out <= 16'hF9EE;    16'd30742: out <= 16'hFDF1;    16'd30743: out <= 16'h06DA;
    16'd30744: out <= 16'hFE4A;    16'd30745: out <= 16'h0127;    16'd30746: out <= 16'h03BF;    16'd30747: out <= 16'h03C9;
    16'd30748: out <= 16'h0035;    16'd30749: out <= 16'h0B7B;    16'd30750: out <= 16'hFD22;    16'd30751: out <= 16'h0172;
    16'd30752: out <= 16'hFB78;    16'd30753: out <= 16'h003F;    16'd30754: out <= 16'h007C;    16'd30755: out <= 16'hFC4A;
    16'd30756: out <= 16'h04E3;    16'd30757: out <= 16'h063D;    16'd30758: out <= 16'hFC22;    16'd30759: out <= 16'hFF2C;
    16'd30760: out <= 16'h043A;    16'd30761: out <= 16'h0367;    16'd30762: out <= 16'h0759;    16'd30763: out <= 16'hFD9C;
    16'd30764: out <= 16'h0877;    16'd30765: out <= 16'h0464;    16'd30766: out <= 16'hFF7B;    16'd30767: out <= 16'h0433;
    16'd30768: out <= 16'h01B3;    16'd30769: out <= 16'h01D8;    16'd30770: out <= 16'h03EB;    16'd30771: out <= 16'h05FC;
    16'd30772: out <= 16'hFDBA;    16'd30773: out <= 16'hFF71;    16'd30774: out <= 16'h05B5;    16'd30775: out <= 16'h0226;
    16'd30776: out <= 16'hFF8F;    16'd30777: out <= 16'h023B;    16'd30778: out <= 16'h03B0;    16'd30779: out <= 16'h05E1;
    16'd30780: out <= 16'h04AA;    16'd30781: out <= 16'h05D5;    16'd30782: out <= 16'h00DC;    16'd30783: out <= 16'hFD87;
    16'd30784: out <= 16'h07E0;    16'd30785: out <= 16'h0313;    16'd30786: out <= 16'hF726;    16'd30787: out <= 16'h0761;
    16'd30788: out <= 16'h0465;    16'd30789: out <= 16'h0175;    16'd30790: out <= 16'h0022;    16'd30791: out <= 16'h0178;
    16'd30792: out <= 16'h0276;    16'd30793: out <= 16'h0BA0;    16'd30794: out <= 16'h08F0;    16'd30795: out <= 16'h04B8;
    16'd30796: out <= 16'h0475;    16'd30797: out <= 16'h0171;    16'd30798: out <= 16'h02A0;    16'd30799: out <= 16'h070D;
    16'd30800: out <= 16'h0842;    16'd30801: out <= 16'h028B;    16'd30802: out <= 16'hFFD0;    16'd30803: out <= 16'h031A;
    16'd30804: out <= 16'hFF9B;    16'd30805: out <= 16'h017F;    16'd30806: out <= 16'h0517;    16'd30807: out <= 16'h06C1;
    16'd30808: out <= 16'h0A39;    16'd30809: out <= 16'h0981;    16'd30810: out <= 16'h022C;    16'd30811: out <= 16'hFFC6;
    16'd30812: out <= 16'hFF2E;    16'd30813: out <= 16'h0413;    16'd30814: out <= 16'h0207;    16'd30815: out <= 16'h0408;
    16'd30816: out <= 16'h042D;    16'd30817: out <= 16'h0605;    16'd30818: out <= 16'h037E;    16'd30819: out <= 16'h05F2;
    16'd30820: out <= 16'h066C;    16'd30821: out <= 16'h07C7;    16'd30822: out <= 16'h0535;    16'd30823: out <= 16'h0242;
    16'd30824: out <= 16'hFEA4;    16'd30825: out <= 16'hFD86;    16'd30826: out <= 16'h02F7;    16'd30827: out <= 16'h0129;
    16'd30828: out <= 16'h01E2;    16'd30829: out <= 16'h018D;    16'd30830: out <= 16'h020D;    16'd30831: out <= 16'h03FE;
    16'd30832: out <= 16'h0906;    16'd30833: out <= 16'h05CC;    16'd30834: out <= 16'h0212;    16'd30835: out <= 16'h0028;
    16'd30836: out <= 16'hFFBB;    16'd30837: out <= 16'h073B;    16'd30838: out <= 16'h0426;    16'd30839: out <= 16'h0637;
    16'd30840: out <= 16'hFE7E;    16'd30841: out <= 16'hF9C4;    16'd30842: out <= 16'h0013;    16'd30843: out <= 16'h010D;
    16'd30844: out <= 16'h07CD;    16'd30845: out <= 16'h0189;    16'd30846: out <= 16'h0200;    16'd30847: out <= 16'h031F;
    16'd30848: out <= 16'h053C;    16'd30849: out <= 16'h03B9;    16'd30850: out <= 16'h0F8F;    16'd30851: out <= 16'h0094;
    16'd30852: out <= 16'hFD63;    16'd30853: out <= 16'h0403;    16'd30854: out <= 16'h0E54;    16'd30855: out <= 16'h0252;
    16'd30856: out <= 16'hFBA0;    16'd30857: out <= 16'h0752;    16'd30858: out <= 16'h03B8;    16'd30859: out <= 16'h05D7;
    16'd30860: out <= 16'h02B0;    16'd30861: out <= 16'h06F5;    16'd30862: out <= 16'h005C;    16'd30863: out <= 16'hFE83;
    16'd30864: out <= 16'h07ED;    16'd30865: out <= 16'h0283;    16'd30866: out <= 16'hFF8A;    16'd30867: out <= 16'h06A1;
    16'd30868: out <= 16'h0463;    16'd30869: out <= 16'h0601;    16'd30870: out <= 16'h02FB;    16'd30871: out <= 16'h025B;
    16'd30872: out <= 16'h0958;    16'd30873: out <= 16'h09B5;    16'd30874: out <= 16'h044F;    16'd30875: out <= 16'h0A1C;
    16'd30876: out <= 16'h0890;    16'd30877: out <= 16'hFDD2;    16'd30878: out <= 16'h053E;    16'd30879: out <= 16'h011D;
    16'd30880: out <= 16'h075E;    16'd30881: out <= 16'h046F;    16'd30882: out <= 16'h092D;    16'd30883: out <= 16'h083E;
    16'd30884: out <= 16'h03DB;    16'd30885: out <= 16'h0405;    16'd30886: out <= 16'h0447;    16'd30887: out <= 16'h028C;
    16'd30888: out <= 16'hFDDC;    16'd30889: out <= 16'h0B01;    16'd30890: out <= 16'h07D4;    16'd30891: out <= 16'h0328;
    16'd30892: out <= 16'hFEB0;    16'd30893: out <= 16'h01EF;    16'd30894: out <= 16'h084A;    16'd30895: out <= 16'h09F4;
    16'd30896: out <= 16'h0BEB;    16'd30897: out <= 16'h0552;    16'd30898: out <= 16'h045B;    16'd30899: out <= 16'h0229;
    16'd30900: out <= 16'h04B6;    16'd30901: out <= 16'h062A;    16'd30902: out <= 16'hFC79;    16'd30903: out <= 16'h07BC;
    16'd30904: out <= 16'h049D;    16'd30905: out <= 16'h0211;    16'd30906: out <= 16'h05D8;    16'd30907: out <= 16'h0BC2;
    16'd30908: out <= 16'h0765;    16'd30909: out <= 16'hFE7F;    16'd30910: out <= 16'h0152;    16'd30911: out <= 16'h017A;
    16'd30912: out <= 16'h0648;    16'd30913: out <= 16'h037C;    16'd30914: out <= 16'hFDDB;    16'd30915: out <= 16'h0414;
    16'd30916: out <= 16'h01C2;    16'd30917: out <= 16'h04A1;    16'd30918: out <= 16'h04B6;    16'd30919: out <= 16'h0912;
    16'd30920: out <= 16'h05CE;    16'd30921: out <= 16'h087D;    16'd30922: out <= 16'hFE24;    16'd30923: out <= 16'hFD05;
    16'd30924: out <= 16'h07F2;    16'd30925: out <= 16'h01C2;    16'd30926: out <= 16'h055D;    16'd30927: out <= 16'h056A;
    16'd30928: out <= 16'hFF3B;    16'd30929: out <= 16'h05B6;    16'd30930: out <= 16'h04C4;    16'd30931: out <= 16'hFABA;
    16'd30932: out <= 16'h0BAE;    16'd30933: out <= 16'h0B6F;    16'd30934: out <= 16'h0504;    16'd30935: out <= 16'h0027;
    16'd30936: out <= 16'hF687;    16'd30937: out <= 16'hFD5B;    16'd30938: out <= 16'h0139;    16'd30939: out <= 16'hF823;
    16'd30940: out <= 16'hFD7B;    16'd30941: out <= 16'h0178;    16'd30942: out <= 16'h004C;    16'd30943: out <= 16'hFF15;
    16'd30944: out <= 16'hF968;    16'd30945: out <= 16'hFC40;    16'd30946: out <= 16'h05A4;    16'd30947: out <= 16'h044C;
    16'd30948: out <= 16'h053F;    16'd30949: out <= 16'h0016;    16'd30950: out <= 16'hFB5B;    16'd30951: out <= 16'h06CC;
    16'd30952: out <= 16'h0691;    16'd30953: out <= 16'h0013;    16'd30954: out <= 16'h05C3;    16'd30955: out <= 16'hFC0E;
    16'd30956: out <= 16'h0344;    16'd30957: out <= 16'h047C;    16'd30958: out <= 16'h0621;    16'd30959: out <= 16'h05B0;
    16'd30960: out <= 16'h057C;    16'd30961: out <= 16'h04AD;    16'd30962: out <= 16'hFFF5;    16'd30963: out <= 16'hFBAC;
    16'd30964: out <= 16'hFEF2;    16'd30965: out <= 16'h0384;    16'd30966: out <= 16'hFDD5;    16'd30967: out <= 16'hFFEA;
    16'd30968: out <= 16'h0044;    16'd30969: out <= 16'hFC5D;    16'd30970: out <= 16'h068C;    16'd30971: out <= 16'h0076;
    16'd30972: out <= 16'h018A;    16'd30973: out <= 16'h031D;    16'd30974: out <= 16'h015E;    16'd30975: out <= 16'hFF90;
    16'd30976: out <= 16'hF4A5;    16'd30977: out <= 16'hFA7F;    16'd30978: out <= 16'hFF4E;    16'd30979: out <= 16'hFC69;
    16'd30980: out <= 16'h012C;    16'd30981: out <= 16'h0048;    16'd30982: out <= 16'h00EA;    16'd30983: out <= 16'h00DB;
    16'd30984: out <= 16'hFDE7;    16'd30985: out <= 16'hFF86;    16'd30986: out <= 16'h0044;    16'd30987: out <= 16'hFF98;
    16'd30988: out <= 16'hFE4E;    16'd30989: out <= 16'hFBE9;    16'd30990: out <= 16'hFFB0;    16'd30991: out <= 16'h0003;
    16'd30992: out <= 16'h0468;    16'd30993: out <= 16'hFCD2;    16'd30994: out <= 16'hFF3A;    16'd30995: out <= 16'h0453;
    16'd30996: out <= 16'h0020;    16'd30997: out <= 16'h06BF;    16'd30998: out <= 16'h0300;    16'd30999: out <= 16'hFDEC;
    16'd31000: out <= 16'hFF17;    16'd31001: out <= 16'h011E;    16'd31002: out <= 16'h0642;    16'd31003: out <= 16'h0313;
    16'd31004: out <= 16'hFD95;    16'd31005: out <= 16'h0522;    16'd31006: out <= 16'hFEB8;    16'd31007: out <= 16'hFF89;
    16'd31008: out <= 16'h0472;    16'd31009: out <= 16'h0723;    16'd31010: out <= 16'h00D8;    16'd31011: out <= 16'h02F7;
    16'd31012: out <= 16'h0542;    16'd31013: out <= 16'h01CA;    16'd31014: out <= 16'hFDC2;    16'd31015: out <= 16'h08DC;
    16'd31016: out <= 16'h01D0;    16'd31017: out <= 16'h0729;    16'd31018: out <= 16'hFDFE;    16'd31019: out <= 16'hFBA6;
    16'd31020: out <= 16'h0444;    16'd31021: out <= 16'h076B;    16'd31022: out <= 16'hFC45;    16'd31023: out <= 16'hFD32;
    16'd31024: out <= 16'h0367;    16'd31025: out <= 16'h03F1;    16'd31026: out <= 16'h02BD;    16'd31027: out <= 16'h0381;
    16'd31028: out <= 16'h01DC;    16'd31029: out <= 16'h0555;    16'd31030: out <= 16'hFFAF;    16'd31031: out <= 16'h0841;
    16'd31032: out <= 16'h0498;    16'd31033: out <= 16'h0BFD;    16'd31034: out <= 16'h0031;    16'd31035: out <= 16'h02C8;
    16'd31036: out <= 16'h0510;    16'd31037: out <= 16'h0099;    16'd31038: out <= 16'hFDF2;    16'd31039: out <= 16'h0700;
    16'd31040: out <= 16'h0FAB;    16'd31041: out <= 16'h07EB;    16'd31042: out <= 16'h07BE;    16'd31043: out <= 16'h00F2;
    16'd31044: out <= 16'h03AB;    16'd31045: out <= 16'h03A1;    16'd31046: out <= 16'h0623;    16'd31047: out <= 16'h0074;
    16'd31048: out <= 16'h033A;    16'd31049: out <= 16'h03A3;    16'd31050: out <= 16'h08CF;    16'd31051: out <= 16'h0281;
    16'd31052: out <= 16'h0672;    16'd31053: out <= 16'h007B;    16'd31054: out <= 16'h03A4;    16'd31055: out <= 16'h04DE;
    16'd31056: out <= 16'h0956;    16'd31057: out <= 16'h0496;    16'd31058: out <= 16'h0A78;    16'd31059: out <= 16'h00A3;
    16'd31060: out <= 16'h06B0;    16'd31061: out <= 16'h09B7;    16'd31062: out <= 16'h00A1;    16'd31063: out <= 16'h0787;
    16'd31064: out <= 16'h052D;    16'd31065: out <= 16'h0353;    16'd31066: out <= 16'h03CE;    16'd31067: out <= 16'h0634;
    16'd31068: out <= 16'h04D8;    16'd31069: out <= 16'h06CC;    16'd31070: out <= 16'h0797;    16'd31071: out <= 16'h0705;
    16'd31072: out <= 16'h0C5A;    16'd31073: out <= 16'h0533;    16'd31074: out <= 16'h02B8;    16'd31075: out <= 16'hFF12;
    16'd31076: out <= 16'hFE7D;    16'd31077: out <= 16'hFF7B;    16'd31078: out <= 16'h07B7;    16'd31079: out <= 16'h032E;
    16'd31080: out <= 16'h066B;    16'd31081: out <= 16'h00B4;    16'd31082: out <= 16'hFE3A;    16'd31083: out <= 16'h0451;
    16'd31084: out <= 16'h076D;    16'd31085: out <= 16'h0263;    16'd31086: out <= 16'hFD67;    16'd31087: out <= 16'h05E7;
    16'd31088: out <= 16'h0326;    16'd31089: out <= 16'h0B3E;    16'd31090: out <= 16'h0216;    16'd31091: out <= 16'hFFCE;
    16'd31092: out <= 16'h0023;    16'd31093: out <= 16'h078F;    16'd31094: out <= 16'h0574;    16'd31095: out <= 16'h0657;
    16'd31096: out <= 16'hFD15;    16'd31097: out <= 16'h0BAC;    16'd31098: out <= 16'h0142;    16'd31099: out <= 16'hFB22;
    16'd31100: out <= 16'h00A0;    16'd31101: out <= 16'h0502;    16'd31102: out <= 16'h076B;    16'd31103: out <= 16'h00A1;
    16'd31104: out <= 16'h07CC;    16'd31105: out <= 16'h02B2;    16'd31106: out <= 16'h0299;    16'd31107: out <= 16'h02D4;
    16'd31108: out <= 16'h081F;    16'd31109: out <= 16'h08A7;    16'd31110: out <= 16'h01AE;    16'd31111: out <= 16'h0562;
    16'd31112: out <= 16'h0430;    16'd31113: out <= 16'h0235;    16'd31114: out <= 16'hFAC6;    16'd31115: out <= 16'h0535;
    16'd31116: out <= 16'h091B;    16'd31117: out <= 16'h00DC;    16'd31118: out <= 16'h0A7F;    16'd31119: out <= 16'hFFCE;
    16'd31120: out <= 16'h0A10;    16'd31121: out <= 16'h0A8C;    16'd31122: out <= 16'h041F;    16'd31123: out <= 16'h0476;
    16'd31124: out <= 16'h0659;    16'd31125: out <= 16'h098F;    16'd31126: out <= 16'h0576;    16'd31127: out <= 16'hFE7A;
    16'd31128: out <= 16'h05C3;    16'd31129: out <= 16'hFCF8;    16'd31130: out <= 16'h0256;    16'd31131: out <= 16'hFBC0;
    16'd31132: out <= 16'h0798;    16'd31133: out <= 16'h03D2;    16'd31134: out <= 16'h0660;    16'd31135: out <= 16'h078B;
    16'd31136: out <= 16'h06BD;    16'd31137: out <= 16'h04BF;    16'd31138: out <= 16'h04FF;    16'd31139: out <= 16'h0467;
    16'd31140: out <= 16'h065A;    16'd31141: out <= 16'h0468;    16'd31142: out <= 16'h0123;    16'd31143: out <= 16'h0A6A;
    16'd31144: out <= 16'h0371;    16'd31145: out <= 16'h0175;    16'd31146: out <= 16'hFF10;    16'd31147: out <= 16'h084B;
    16'd31148: out <= 16'h09B0;    16'd31149: out <= 16'h0701;    16'd31150: out <= 16'h059D;    16'd31151: out <= 16'h0379;
    16'd31152: out <= 16'h0645;    16'd31153: out <= 16'h0792;    16'd31154: out <= 16'h04E3;    16'd31155: out <= 16'h0493;
    16'd31156: out <= 16'hFCC1;    16'd31157: out <= 16'hFFEB;    16'd31158: out <= 16'h0523;    16'd31159: out <= 16'h03DB;
    16'd31160: out <= 16'h01F2;    16'd31161: out <= 16'h0A3C;    16'd31162: out <= 16'h029A;    16'd31163: out <= 16'h06A0;
    16'd31164: out <= 16'h00DB;    16'd31165: out <= 16'h06C4;    16'd31166: out <= 16'h017B;    16'd31167: out <= 16'h00BA;
    16'd31168: out <= 16'h07A8;    16'd31169: out <= 16'h02EF;    16'd31170: out <= 16'h0120;    16'd31171: out <= 16'h0A6C;
    16'd31172: out <= 16'h0090;    16'd31173: out <= 16'h01D4;    16'd31174: out <= 16'h0517;    16'd31175: out <= 16'h0680;
    16'd31176: out <= 16'h0656;    16'd31177: out <= 16'h00A3;    16'd31178: out <= 16'hFDCB;    16'd31179: out <= 16'h024F;
    16'd31180: out <= 16'h0222;    16'd31181: out <= 16'h0773;    16'd31182: out <= 16'h0756;    16'd31183: out <= 16'h0317;
    16'd31184: out <= 16'h0417;    16'd31185: out <= 16'h0043;    16'd31186: out <= 16'h04DF;    16'd31187: out <= 16'hFDAB;
    16'd31188: out <= 16'h0341;    16'd31189: out <= 16'h0682;    16'd31190: out <= 16'h02C0;    16'd31191: out <= 16'h0444;
    16'd31192: out <= 16'h06BF;    16'd31193: out <= 16'h01E0;    16'd31194: out <= 16'h0219;    16'd31195: out <= 16'hFFC4;
    16'd31196: out <= 16'hFBC0;    16'd31197: out <= 16'hFA25;    16'd31198: out <= 16'hFC09;    16'd31199: out <= 16'h0157;
    16'd31200: out <= 16'hFFFE;    16'd31201: out <= 16'h01AB;    16'd31202: out <= 16'h00F0;    16'd31203: out <= 16'hFF8A;
    16'd31204: out <= 16'hFF98;    16'd31205: out <= 16'h095B;    16'd31206: out <= 16'h0A31;    16'd31207: out <= 16'h04FE;
    16'd31208: out <= 16'hFC1D;    16'd31209: out <= 16'hF6F9;    16'd31210: out <= 16'hF8AE;    16'd31211: out <= 16'h072B;
    16'd31212: out <= 16'h0672;    16'd31213: out <= 16'hF66C;    16'd31214: out <= 16'h009F;    16'd31215: out <= 16'hFCEA;
    16'd31216: out <= 16'hFC86;    16'd31217: out <= 16'h089A;    16'd31218: out <= 16'hF6E6;    16'd31219: out <= 16'h0252;
    16'd31220: out <= 16'hF8DB;    16'd31221: out <= 16'hFC55;    16'd31222: out <= 16'hFEEB;    16'd31223: out <= 16'hFC84;
    16'd31224: out <= 16'hFD88;    16'd31225: out <= 16'hFF1E;    16'd31226: out <= 16'hFD3E;    16'd31227: out <= 16'hFF0C;
    16'd31228: out <= 16'h0320;    16'd31229: out <= 16'h06DC;    16'd31230: out <= 16'h059D;    16'd31231: out <= 16'hFF71;
    16'd31232: out <= 16'hFBC5;    16'd31233: out <= 16'h0672;    16'd31234: out <= 16'h0461;    16'd31235: out <= 16'hFCDA;
    16'd31236: out <= 16'hFE03;    16'd31237: out <= 16'hFAB3;    16'd31238: out <= 16'h01DD;    16'd31239: out <= 16'h028F;
    16'd31240: out <= 16'h06F7;    16'd31241: out <= 16'hFCBD;    16'd31242: out <= 16'hFF09;    16'd31243: out <= 16'hFE47;
    16'd31244: out <= 16'h0932;    16'd31245: out <= 16'h008B;    16'd31246: out <= 16'hFF09;    16'd31247: out <= 16'h000C;
    16'd31248: out <= 16'h0032;    16'd31249: out <= 16'hFEF2;    16'd31250: out <= 16'h0374;    16'd31251: out <= 16'hF8C3;
    16'd31252: out <= 16'hF757;    16'd31253: out <= 16'h01E7;    16'd31254: out <= 16'h010B;    16'd31255: out <= 16'h065A;
    16'd31256: out <= 16'h0042;    16'd31257: out <= 16'h039A;    16'd31258: out <= 16'h002F;    16'd31259: out <= 16'hFD37;
    16'd31260: out <= 16'hFCB3;    16'd31261: out <= 16'h07BB;    16'd31262: out <= 16'h00DE;    16'd31263: out <= 16'h06AC;
    16'd31264: out <= 16'h03C0;    16'd31265: out <= 16'h0162;    16'd31266: out <= 16'h04E5;    16'd31267: out <= 16'h0741;
    16'd31268: out <= 16'h08BC;    16'd31269: out <= 16'h0460;    16'd31270: out <= 16'h03A9;    16'd31271: out <= 16'h02D1;
    16'd31272: out <= 16'h074A;    16'd31273: out <= 16'h04AE;    16'd31274: out <= 16'h0522;    16'd31275: out <= 16'h0277;
    16'd31276: out <= 16'h056F;    16'd31277: out <= 16'h0309;    16'd31278: out <= 16'h027E;    16'd31279: out <= 16'h084F;
    16'd31280: out <= 16'hFD18;    16'd31281: out <= 16'h0376;    16'd31282: out <= 16'h002F;    16'd31283: out <= 16'h0379;
    16'd31284: out <= 16'hFB01;    16'd31285: out <= 16'hFEE3;    16'd31286: out <= 16'hF72A;    16'd31287: out <= 16'h024B;
    16'd31288: out <= 16'h073E;    16'd31289: out <= 16'h0B7C;    16'd31290: out <= 16'h06A2;    16'd31291: out <= 16'h02D1;
    16'd31292: out <= 16'h020F;    16'd31293: out <= 16'h0746;    16'd31294: out <= 16'h0064;    16'd31295: out <= 16'hFF4B;
    16'd31296: out <= 16'h0238;    16'd31297: out <= 16'h015D;    16'd31298: out <= 16'h085A;    16'd31299: out <= 16'h049D;
    16'd31300: out <= 16'h01B1;    16'd31301: out <= 16'hFE2C;    16'd31302: out <= 16'h02C3;    16'd31303: out <= 16'hFB77;
    16'd31304: out <= 16'h0444;    16'd31305: out <= 16'h0172;    16'd31306: out <= 16'h011F;    16'd31307: out <= 16'h01C8;
    16'd31308: out <= 16'h0AEE;    16'd31309: out <= 16'h03CF;    16'd31310: out <= 16'hFF5A;    16'd31311: out <= 16'h055D;
    16'd31312: out <= 16'h054E;    16'd31313: out <= 16'h0474;    16'd31314: out <= 16'hFEB3;    16'd31315: out <= 16'h03EA;
    16'd31316: out <= 16'h05C9;    16'd31317: out <= 16'h00FC;    16'd31318: out <= 16'h035D;    16'd31319: out <= 16'h05BD;
    16'd31320: out <= 16'hFE16;    16'd31321: out <= 16'h00B2;    16'd31322: out <= 16'hFD4B;    16'd31323: out <= 16'h02C2;
    16'd31324: out <= 16'h0504;    16'd31325: out <= 16'h08EB;    16'd31326: out <= 16'h0780;    16'd31327: out <= 16'h04B7;
    16'd31328: out <= 16'h0504;    16'd31329: out <= 16'h0165;    16'd31330: out <= 16'h0579;    16'd31331: out <= 16'hFE12;
    16'd31332: out <= 16'h0377;    16'd31333: out <= 16'h0907;    16'd31334: out <= 16'hFC3F;    16'd31335: out <= 16'hFF80;
    16'd31336: out <= 16'h042E;    16'd31337: out <= 16'h0AFB;    16'd31338: out <= 16'h0836;    16'd31339: out <= 16'h05E3;
    16'd31340: out <= 16'h00AD;    16'd31341: out <= 16'h0601;    16'd31342: out <= 16'h0819;    16'd31343: out <= 16'h0950;
    16'd31344: out <= 16'h00D7;    16'd31345: out <= 16'h036A;    16'd31346: out <= 16'hFF1F;    16'd31347: out <= 16'h0353;
    16'd31348: out <= 16'h02BC;    16'd31349: out <= 16'h0136;    16'd31350: out <= 16'h02C8;    16'd31351: out <= 16'h051E;
    16'd31352: out <= 16'h003A;    16'd31353: out <= 16'h01A1;    16'd31354: out <= 16'h056B;    16'd31355: out <= 16'h076D;
    16'd31356: out <= 16'hFCF3;    16'd31357: out <= 16'hFFDF;    16'd31358: out <= 16'hFD1E;    16'd31359: out <= 16'h02D2;
    16'd31360: out <= 16'h0185;    16'd31361: out <= 16'h0047;    16'd31362: out <= 16'h0210;    16'd31363: out <= 16'h05AA;
    16'd31364: out <= 16'hFF09;    16'd31365: out <= 16'h011B;    16'd31366: out <= 16'h036D;    16'd31367: out <= 16'h035D;
    16'd31368: out <= 16'h06CA;    16'd31369: out <= 16'h0265;    16'd31370: out <= 16'hFDC9;    16'd31371: out <= 16'h0508;
    16'd31372: out <= 16'h041F;    16'd31373: out <= 16'h057B;    16'd31374: out <= 16'h0691;    16'd31375: out <= 16'h0B6B;
    16'd31376: out <= 16'hFED4;    16'd31377: out <= 16'h03D1;    16'd31378: out <= 16'h0574;    16'd31379: out <= 16'h030C;
    16'd31380: out <= 16'hFD8D;    16'd31381: out <= 16'h0295;    16'd31382: out <= 16'h0A70;    16'd31383: out <= 16'h0182;
    16'd31384: out <= 16'h0922;    16'd31385: out <= 16'h0434;    16'd31386: out <= 16'h01CE;    16'd31387: out <= 16'h07E0;
    16'd31388: out <= 16'h0760;    16'd31389: out <= 16'h0641;    16'd31390: out <= 16'h0C2A;    16'd31391: out <= 16'h01D4;
    16'd31392: out <= 16'h042C;    16'd31393: out <= 16'hFE53;    16'd31394: out <= 16'h031C;    16'd31395: out <= 16'h0018;
    16'd31396: out <= 16'h01A6;    16'd31397: out <= 16'hFE5F;    16'd31398: out <= 16'h0574;    16'd31399: out <= 16'h049B;
    16'd31400: out <= 16'h05D3;    16'd31401: out <= 16'h0579;    16'd31402: out <= 16'h048B;    16'd31403: out <= 16'h04FC;
    16'd31404: out <= 16'hFFD2;    16'd31405: out <= 16'h0834;    16'd31406: out <= 16'h00C1;    16'd31407: out <= 16'h0AB4;
    16'd31408: out <= 16'h0028;    16'd31409: out <= 16'h0234;    16'd31410: out <= 16'h06DE;    16'd31411: out <= 16'hFCF3;
    16'd31412: out <= 16'hFED5;    16'd31413: out <= 16'h0422;    16'd31414: out <= 16'hFFD9;    16'd31415: out <= 16'h056B;
    16'd31416: out <= 16'h042A;    16'd31417: out <= 16'h0A25;    16'd31418: out <= 16'hFD3D;    16'd31419: out <= 16'h089E;
    16'd31420: out <= 16'h0696;    16'd31421: out <= 16'hFFFD;    16'd31422: out <= 16'h0BC6;    16'd31423: out <= 16'hFF19;
    16'd31424: out <= 16'h05E0;    16'd31425: out <= 16'h0570;    16'd31426: out <= 16'h0297;    16'd31427: out <= 16'h085B;
    16'd31428: out <= 16'h064E;    16'd31429: out <= 16'h03E3;    16'd31430: out <= 16'h08EE;    16'd31431: out <= 16'h0AC8;
    16'd31432: out <= 16'h0323;    16'd31433: out <= 16'h0474;    16'd31434: out <= 16'h031E;    16'd31435: out <= 16'h0759;
    16'd31436: out <= 16'hFCBA;    16'd31437: out <= 16'h08A5;    16'd31438: out <= 16'h02D2;    16'd31439: out <= 16'h014F;
    16'd31440: out <= 16'h02A4;    16'd31441: out <= 16'hFBE8;    16'd31442: out <= 16'h0704;    16'd31443: out <= 16'h04A0;
    16'd31444: out <= 16'h02B2;    16'd31445: out <= 16'h025D;    16'd31446: out <= 16'hFC84;    16'd31447: out <= 16'hFDE1;
    16'd31448: out <= 16'hFC90;    16'd31449: out <= 16'h01A2;    16'd31450: out <= 16'hFE03;    16'd31451: out <= 16'h06EC;
    16'd31452: out <= 16'h066E;    16'd31453: out <= 16'h0270;    16'd31454: out <= 16'h04D1;    16'd31455: out <= 16'h055B;
    16'd31456: out <= 16'h03AC;    16'd31457: out <= 16'h06AF;    16'd31458: out <= 16'h055B;    16'd31459: out <= 16'h082E;
    16'd31460: out <= 16'h0164;    16'd31461: out <= 16'h0020;    16'd31462: out <= 16'h05C5;    16'd31463: out <= 16'h026D;
    16'd31464: out <= 16'hFF2F;    16'd31465: out <= 16'h062D;    16'd31466: out <= 16'h023B;    16'd31467: out <= 16'hFDFB;
    16'd31468: out <= 16'h03A8;    16'd31469: out <= 16'h0150;    16'd31470: out <= 16'h04A8;    16'd31471: out <= 16'h0286;
    16'd31472: out <= 16'h01E3;    16'd31473: out <= 16'h00E8;    16'd31474: out <= 16'hF95C;    16'd31475: out <= 16'h03B4;
    16'd31476: out <= 16'h01E3;    16'd31477: out <= 16'h03BB;    16'd31478: out <= 16'h0566;    16'd31479: out <= 16'hF928;
    16'd31480: out <= 16'h053A;    16'd31481: out <= 16'h03AC;    16'd31482: out <= 16'hFF54;    16'd31483: out <= 16'h01D5;
    16'd31484: out <= 16'hFADB;    16'd31485: out <= 16'hF5EF;    16'd31486: out <= 16'h010C;    16'd31487: out <= 16'h0238;
    16'd31488: out <= 16'h021A;    16'd31489: out <= 16'hFC05;    16'd31490: out <= 16'hFE49;    16'd31491: out <= 16'hFB9D;
    16'd31492: out <= 16'hFFBC;    16'd31493: out <= 16'h0207;    16'd31494: out <= 16'h0150;    16'd31495: out <= 16'hFF01;
    16'd31496: out <= 16'hFE58;    16'd31497: out <= 16'h06A3;    16'd31498: out <= 16'h0213;    16'd31499: out <= 16'hFE71;
    16'd31500: out <= 16'h077B;    16'd31501: out <= 16'h0172;    16'd31502: out <= 16'h050B;    16'd31503: out <= 16'hFF1F;
    16'd31504: out <= 16'hFE07;    16'd31505: out <= 16'h0289;    16'd31506: out <= 16'hFC13;    16'd31507: out <= 16'h0659;
    16'd31508: out <= 16'h0862;    16'd31509: out <= 16'h0122;    16'd31510: out <= 16'h003E;    16'd31511: out <= 16'h0769;
    16'd31512: out <= 16'hFF2C;    16'd31513: out <= 16'h0379;    16'd31514: out <= 16'h01EF;    16'd31515: out <= 16'h0357;
    16'd31516: out <= 16'h025E;    16'd31517: out <= 16'h0574;    16'd31518: out <= 16'h0833;    16'd31519: out <= 16'h070F;
    16'd31520: out <= 16'h0880;    16'd31521: out <= 16'hFEE9;    16'd31522: out <= 16'h03C3;    16'd31523: out <= 16'hFE0E;
    16'd31524: out <= 16'h05D0;    16'd31525: out <= 16'h0427;    16'd31526: out <= 16'h0DA5;    16'd31527: out <= 16'h089E;
    16'd31528: out <= 16'h0909;    16'd31529: out <= 16'h0127;    16'd31530: out <= 16'h043F;    16'd31531: out <= 16'h06F7;
    16'd31532: out <= 16'hFEDF;    16'd31533: out <= 16'h0AE2;    16'd31534: out <= 16'h0580;    16'd31535: out <= 16'hFE6D;
    16'd31536: out <= 16'h046D;    16'd31537: out <= 16'h0827;    16'd31538: out <= 16'h046F;    16'd31539: out <= 16'h0250;
    16'd31540: out <= 16'h078D;    16'd31541: out <= 16'h05A1;    16'd31542: out <= 16'h06EF;    16'd31543: out <= 16'h0EFB;
    16'd31544: out <= 16'h066F;    16'd31545: out <= 16'h051F;    16'd31546: out <= 16'h07E9;    16'd31547: out <= 16'h0653;
    16'd31548: out <= 16'h0695;    16'd31549: out <= 16'h063D;    16'd31550: out <= 16'hFAB0;    16'd31551: out <= 16'h0152;
    16'd31552: out <= 16'h0463;    16'd31553: out <= 16'h03BF;    16'd31554: out <= 16'h02A2;    16'd31555: out <= 16'h008D;
    16'd31556: out <= 16'hFD79;    16'd31557: out <= 16'h03E5;    16'd31558: out <= 16'h03AB;    16'd31559: out <= 16'hFFA7;
    16'd31560: out <= 16'hFA5D;    16'd31561: out <= 16'h01F6;    16'd31562: out <= 16'h0502;    16'd31563: out <= 16'hFD34;
    16'd31564: out <= 16'h06D4;    16'd31565: out <= 16'h0052;    16'd31566: out <= 16'h0C5E;    16'd31567: out <= 16'h08AE;
    16'd31568: out <= 16'h0597;    16'd31569: out <= 16'hFE5B;    16'd31570: out <= 16'h0843;    16'd31571: out <= 16'h08FA;
    16'd31572: out <= 16'hFFE8;    16'd31573: out <= 16'h0AB2;    16'd31574: out <= 16'h0725;    16'd31575: out <= 16'h0640;
    16'd31576: out <= 16'h0399;    16'd31577: out <= 16'h03F4;    16'd31578: out <= 16'hF9D6;    16'd31579: out <= 16'h077A;
    16'd31580: out <= 16'hFD4A;    16'd31581: out <= 16'hFE36;    16'd31582: out <= 16'h020B;    16'd31583: out <= 16'h0211;
    16'd31584: out <= 16'h0528;    16'd31585: out <= 16'h028C;    16'd31586: out <= 16'h0463;    16'd31587: out <= 16'h05E2;
    16'd31588: out <= 16'h050B;    16'd31589: out <= 16'h0018;    16'd31590: out <= 16'h0B2D;    16'd31591: out <= 16'h0656;
    16'd31592: out <= 16'hFEA7;    16'd31593: out <= 16'h04D5;    16'd31594: out <= 16'h021A;    16'd31595: out <= 16'hFFF5;
    16'd31596: out <= 16'h0239;    16'd31597: out <= 16'hFB91;    16'd31598: out <= 16'h02B3;    16'd31599: out <= 16'h0765;
    16'd31600: out <= 16'h077F;    16'd31601: out <= 16'h0509;    16'd31602: out <= 16'h00BB;    16'd31603: out <= 16'h0444;
    16'd31604: out <= 16'h0234;    16'd31605: out <= 16'h050E;    16'd31606: out <= 16'h066E;    16'd31607: out <= 16'h0063;
    16'd31608: out <= 16'h0C99;    16'd31609: out <= 16'hFA8F;    16'd31610: out <= 16'hFDD6;    16'd31611: out <= 16'h0A0C;
    16'd31612: out <= 16'hFC22;    16'd31613: out <= 16'h06C6;    16'd31614: out <= 16'h06B4;    16'd31615: out <= 16'h045A;
    16'd31616: out <= 16'h0574;    16'd31617: out <= 16'h0016;    16'd31618: out <= 16'h0553;    16'd31619: out <= 16'h0948;
    16'd31620: out <= 16'hFCF2;    16'd31621: out <= 16'h06BC;    16'd31622: out <= 16'h065C;    16'd31623: out <= 16'hFF92;
    16'd31624: out <= 16'h0C2E;    16'd31625: out <= 16'h06E3;    16'd31626: out <= 16'h0277;    16'd31627: out <= 16'h08BE;
    16'd31628: out <= 16'h05E8;    16'd31629: out <= 16'h09D7;    16'd31630: out <= 16'h069C;    16'd31631: out <= 16'h0753;
    16'd31632: out <= 16'h0A1B;    16'd31633: out <= 16'h0101;    16'd31634: out <= 16'h0356;    16'd31635: out <= 16'h03F2;
    16'd31636: out <= 16'h06DE;    16'd31637: out <= 16'h061E;    16'd31638: out <= 16'h0341;    16'd31639: out <= 16'h0456;
    16'd31640: out <= 16'h05A8;    16'd31641: out <= 16'h0678;    16'd31642: out <= 16'h05B6;    16'd31643: out <= 16'h087A;
    16'd31644: out <= 16'h02A7;    16'd31645: out <= 16'h02B9;    16'd31646: out <= 16'h051F;    16'd31647: out <= 16'hFEF8;
    16'd31648: out <= 16'h00BF;    16'd31649: out <= 16'h05C6;    16'd31650: out <= 16'h04C3;    16'd31651: out <= 16'h01EA;
    16'd31652: out <= 16'h0413;    16'd31653: out <= 16'h021F;    16'd31654: out <= 16'h0BDE;    16'd31655: out <= 16'h0888;
    16'd31656: out <= 16'h0253;    16'd31657: out <= 16'hFC19;    16'd31658: out <= 16'h04D1;    16'd31659: out <= 16'h049B;
    16'd31660: out <= 16'h06B2;    16'd31661: out <= 16'hFC96;    16'd31662: out <= 16'h0426;    16'd31663: out <= 16'h0743;
    16'd31664: out <= 16'h03E8;    16'd31665: out <= 16'h075F;    16'd31666: out <= 16'h043E;    16'd31667: out <= 16'h0161;
    16'd31668: out <= 16'hFFF9;    16'd31669: out <= 16'h090F;    16'd31670: out <= 16'h0718;    16'd31671: out <= 16'h05D0;
    16'd31672: out <= 16'h013A;    16'd31673: out <= 16'h00B4;    16'd31674: out <= 16'h00C1;    16'd31675: out <= 16'h03D5;
    16'd31676: out <= 16'h0656;    16'd31677: out <= 16'h06EC;    16'd31678: out <= 16'h09A2;    16'd31679: out <= 16'h021F;
    16'd31680: out <= 16'h055C;    16'd31681: out <= 16'hFB6F;    16'd31682: out <= 16'h01FF;    16'd31683: out <= 16'h03F0;
    16'd31684: out <= 16'h051B;    16'd31685: out <= 16'h04FE;    16'd31686: out <= 16'h04FD;    16'd31687: out <= 16'h037A;
    16'd31688: out <= 16'h03AE;    16'd31689: out <= 16'h0AAE;    16'd31690: out <= 16'h01B8;    16'd31691: out <= 16'h070A;
    16'd31692: out <= 16'h020F;    16'd31693: out <= 16'h07FC;    16'd31694: out <= 16'h08BF;    16'd31695: out <= 16'h010C;
    16'd31696: out <= 16'h0197;    16'd31697: out <= 16'h058C;    16'd31698: out <= 16'h0649;    16'd31699: out <= 16'h03B9;
    16'd31700: out <= 16'h03FF;    16'd31701: out <= 16'h0390;    16'd31702: out <= 16'hFD8B;    16'd31703: out <= 16'h04FF;
    16'd31704: out <= 16'h0486;    16'd31705: out <= 16'h068F;    16'd31706: out <= 16'h05F9;    16'd31707: out <= 16'h01DE;
    16'd31708: out <= 16'h05A5;    16'd31709: out <= 16'hFF84;    16'd31710: out <= 16'h0026;    16'd31711: out <= 16'h06AF;
    16'd31712: out <= 16'h028D;    16'd31713: out <= 16'h0077;    16'd31714: out <= 16'h04D7;    16'd31715: out <= 16'h0973;
    16'd31716: out <= 16'h0401;    16'd31717: out <= 16'h0538;    16'd31718: out <= 16'h0017;    16'd31719: out <= 16'hFA7C;
    16'd31720: out <= 16'hF8B1;    16'd31721: out <= 16'hFCCB;    16'd31722: out <= 16'hFE8C;    16'd31723: out <= 16'h02A1;
    16'd31724: out <= 16'h0698;    16'd31725: out <= 16'h02B4;    16'd31726: out <= 16'h0023;    16'd31727: out <= 16'hFEAA;
    16'd31728: out <= 16'h09AC;    16'd31729: out <= 16'h03B4;    16'd31730: out <= 16'h0888;    16'd31731: out <= 16'hFD8D;
    16'd31732: out <= 16'h065D;    16'd31733: out <= 16'hFE96;    16'd31734: out <= 16'hFB11;    16'd31735: out <= 16'h06DE;
    16'd31736: out <= 16'hFF72;    16'd31737: out <= 16'h0328;    16'd31738: out <= 16'hF633;    16'd31739: out <= 16'hFBC1;
    16'd31740: out <= 16'hFFEC;    16'd31741: out <= 16'h03D3;    16'd31742: out <= 16'h01B3;    16'd31743: out <= 16'hFE8F;
    16'd31744: out <= 16'hFD1F;    16'd31745: out <= 16'h0191;    16'd31746: out <= 16'h06B6;    16'd31747: out <= 16'h0332;
    16'd31748: out <= 16'h00BD;    16'd31749: out <= 16'h0567;    16'd31750: out <= 16'h038F;    16'd31751: out <= 16'hF8E4;
    16'd31752: out <= 16'h0097;    16'd31753: out <= 16'hFDC5;    16'd31754: out <= 16'hFE53;    16'd31755: out <= 16'h0112;
    16'd31756: out <= 16'h0357;    16'd31757: out <= 16'h066A;    16'd31758: out <= 16'hFBC9;    16'd31759: out <= 16'hFE77;
    16'd31760: out <= 16'h0065;    16'd31761: out <= 16'h02C4;    16'd31762: out <= 16'h016C;    16'd31763: out <= 16'hFE64;
    16'd31764: out <= 16'h0AC1;    16'd31765: out <= 16'h089C;    16'd31766: out <= 16'hFAAB;    16'd31767: out <= 16'h0883;
    16'd31768: out <= 16'h09B5;    16'd31769: out <= 16'h012E;    16'd31770: out <= 16'h0D25;    16'd31771: out <= 16'h0013;
    16'd31772: out <= 16'h01F5;    16'd31773: out <= 16'hFFAD;    16'd31774: out <= 16'h0179;    16'd31775: out <= 16'h08F0;
    16'd31776: out <= 16'h00AC;    16'd31777: out <= 16'h051E;    16'd31778: out <= 16'h0376;    16'd31779: out <= 16'h01C2;
    16'd31780: out <= 16'h06CE;    16'd31781: out <= 16'h0722;    16'd31782: out <= 16'h0326;    16'd31783: out <= 16'hFFD2;
    16'd31784: out <= 16'h0658;    16'd31785: out <= 16'h01C3;    16'd31786: out <= 16'h026C;    16'd31787: out <= 16'h0511;
    16'd31788: out <= 16'hFC02;    16'd31789: out <= 16'h058C;    16'd31790: out <= 16'h03A4;    16'd31791: out <= 16'h0567;
    16'd31792: out <= 16'h0560;    16'd31793: out <= 16'h023E;    16'd31794: out <= 16'h01F1;    16'd31795: out <= 16'hFF62;
    16'd31796: out <= 16'h0326;    16'd31797: out <= 16'h031B;    16'd31798: out <= 16'hFDDC;    16'd31799: out <= 16'h06E9;
    16'd31800: out <= 16'h0680;    16'd31801: out <= 16'h00AB;    16'd31802: out <= 16'h01FF;    16'd31803: out <= 16'h032B;
    16'd31804: out <= 16'h0487;    16'd31805: out <= 16'h0A91;    16'd31806: out <= 16'h0660;    16'd31807: out <= 16'h00DF;
    16'd31808: out <= 16'h0841;    16'd31809: out <= 16'h04AE;    16'd31810: out <= 16'h0A6E;    16'd31811: out <= 16'h0921;
    16'd31812: out <= 16'h0548;    16'd31813: out <= 16'hFFBC;    16'd31814: out <= 16'h0158;    16'd31815: out <= 16'h04BF;
    16'd31816: out <= 16'h0392;    16'd31817: out <= 16'h0411;    16'd31818: out <= 16'h0198;    16'd31819: out <= 16'hF781;
    16'd31820: out <= 16'h0211;    16'd31821: out <= 16'h012E;    16'd31822: out <= 16'h0624;    16'd31823: out <= 16'h032D;
    16'd31824: out <= 16'h0BF1;    16'd31825: out <= 16'h035B;    16'd31826: out <= 16'hFD08;    16'd31827: out <= 16'h0799;
    16'd31828: out <= 16'h027C;    16'd31829: out <= 16'h0482;    16'd31830: out <= 16'h03AB;    16'd31831: out <= 16'h03F9;
    16'd31832: out <= 16'hFEFF;    16'd31833: out <= 16'h0621;    16'd31834: out <= 16'h052A;    16'd31835: out <= 16'h0B94;
    16'd31836: out <= 16'h018B;    16'd31837: out <= 16'h04DA;    16'd31838: out <= 16'h04C2;    16'd31839: out <= 16'h02B4;
    16'd31840: out <= 16'h0606;    16'd31841: out <= 16'h06AD;    16'd31842: out <= 16'hFC14;    16'd31843: out <= 16'h0B1F;
    16'd31844: out <= 16'h048D;    16'd31845: out <= 16'h0257;    16'd31846: out <= 16'h0482;    16'd31847: out <= 16'h026D;
    16'd31848: out <= 16'h086F;    16'd31849: out <= 16'h07EB;    16'd31850: out <= 16'h0314;    16'd31851: out <= 16'h05FC;
    16'd31852: out <= 16'h0168;    16'd31853: out <= 16'h0369;    16'd31854: out <= 16'h02E5;    16'd31855: out <= 16'hFE1F;
    16'd31856: out <= 16'h0288;    16'd31857: out <= 16'h092A;    16'd31858: out <= 16'h0745;    16'd31859: out <= 16'h033A;
    16'd31860: out <= 16'h02A3;    16'd31861: out <= 16'h0032;    16'd31862: out <= 16'hFFC2;    16'd31863: out <= 16'h0021;
    16'd31864: out <= 16'h02F7;    16'd31865: out <= 16'h013E;    16'd31866: out <= 16'h04A4;    16'd31867: out <= 16'h01C1;
    16'd31868: out <= 16'h0290;    16'd31869: out <= 16'h0786;    16'd31870: out <= 16'h0712;    16'd31871: out <= 16'h0119;
    16'd31872: out <= 16'h011F;    16'd31873: out <= 16'h01A9;    16'd31874: out <= 16'hFDCA;    16'd31875: out <= 16'h0483;
    16'd31876: out <= 16'h0B0A;    16'd31877: out <= 16'h02AA;    16'd31878: out <= 16'h082D;    16'd31879: out <= 16'h02A4;
    16'd31880: out <= 16'h0BD0;    16'd31881: out <= 16'hFF8F;    16'd31882: out <= 16'h09D2;    16'd31883: out <= 16'h0307;
    16'd31884: out <= 16'h09AD;    16'd31885: out <= 16'h0087;    16'd31886: out <= 16'h0314;    16'd31887: out <= 16'h08FB;
    16'd31888: out <= 16'h04E8;    16'd31889: out <= 16'h043A;    16'd31890: out <= 16'hFC8E;    16'd31891: out <= 16'h0124;
    16'd31892: out <= 16'h040E;    16'd31893: out <= 16'h040B;    16'd31894: out <= 16'h090B;    16'd31895: out <= 16'h02D3;
    16'd31896: out <= 16'h012A;    16'd31897: out <= 16'h0025;    16'd31898: out <= 16'h05A4;    16'd31899: out <= 16'h056F;
    16'd31900: out <= 16'h02F4;    16'd31901: out <= 16'h0845;    16'd31902: out <= 16'h0088;    16'd31903: out <= 16'h00F1;
    16'd31904: out <= 16'h050F;    16'd31905: out <= 16'h0540;    16'd31906: out <= 16'hFEFF;    16'd31907: out <= 16'h0399;
    16'd31908: out <= 16'h0598;    16'd31909: out <= 16'hFE9D;    16'd31910: out <= 16'h0065;    16'd31911: out <= 16'h0771;
    16'd31912: out <= 16'h0086;    16'd31913: out <= 16'h0575;    16'd31914: out <= 16'h0303;    16'd31915: out <= 16'h0681;
    16'd31916: out <= 16'h0451;    16'd31917: out <= 16'h06A2;    16'd31918: out <= 16'h05C0;    16'd31919: out <= 16'hFF83;
    16'd31920: out <= 16'hFFAD;    16'd31921: out <= 16'h00A3;    16'd31922: out <= 16'h054D;    16'd31923: out <= 16'h031F;
    16'd31924: out <= 16'h04D1;    16'd31925: out <= 16'h079A;    16'd31926: out <= 16'h02D2;    16'd31927: out <= 16'h0120;
    16'd31928: out <= 16'h011F;    16'd31929: out <= 16'h098E;    16'd31930: out <= 16'h0343;    16'd31931: out <= 16'h0297;
    16'd31932: out <= 16'h04CF;    16'd31933: out <= 16'h0368;    16'd31934: out <= 16'h05D0;    16'd31935: out <= 16'h0254;
    16'd31936: out <= 16'h0480;    16'd31937: out <= 16'h0573;    16'd31938: out <= 16'h01A6;    16'd31939: out <= 16'h023D;
    16'd31940: out <= 16'h03FF;    16'd31941: out <= 16'h0452;    16'd31942: out <= 16'h02AA;    16'd31943: out <= 16'hFAC5;
    16'd31944: out <= 16'h0369;    16'd31945: out <= 16'hFFC4;    16'd31946: out <= 16'hFB40;    16'd31947: out <= 16'h05E7;
    16'd31948: out <= 16'h0883;    16'd31949: out <= 16'hFCCE;    16'd31950: out <= 16'hFC61;    16'd31951: out <= 16'h06A6;
    16'd31952: out <= 16'h035E;    16'd31953: out <= 16'h0238;    16'd31954: out <= 16'h0839;    16'd31955: out <= 16'h0520;
    16'd31956: out <= 16'h0454;    16'd31957: out <= 16'h095E;    16'd31958: out <= 16'h0084;    16'd31959: out <= 16'h0796;
    16'd31960: out <= 16'h0566;    16'd31961: out <= 16'h03D7;    16'd31962: out <= 16'h0348;    16'd31963: out <= 16'hFB20;
    16'd31964: out <= 16'hFCBC;    16'd31965: out <= 16'hFD9B;    16'd31966: out <= 16'h0217;    16'd31967: out <= 16'h050F;
    16'd31968: out <= 16'h074A;    16'd31969: out <= 16'h06D6;    16'd31970: out <= 16'h07C5;    16'd31971: out <= 16'h01B4;
    16'd31972: out <= 16'hFEB2;    16'd31973: out <= 16'h041B;    16'd31974: out <= 16'h0597;    16'd31975: out <= 16'hFE0A;
    16'd31976: out <= 16'h0418;    16'd31977: out <= 16'h020A;    16'd31978: out <= 16'h047C;    16'd31979: out <= 16'h04D6;
    16'd31980: out <= 16'hFF4B;    16'd31981: out <= 16'hFD7C;    16'd31982: out <= 16'hFE5D;    16'd31983: out <= 16'h014D;
    16'd31984: out <= 16'h006D;    16'd31985: out <= 16'hFE37;    16'd31986: out <= 16'hFC85;    16'd31987: out <= 16'h0107;
    16'd31988: out <= 16'hFA40;    16'd31989: out <= 16'h02D1;    16'd31990: out <= 16'h010D;    16'd31991: out <= 16'h06C8;
    16'd31992: out <= 16'h008C;    16'd31993: out <= 16'hFF21;    16'd31994: out <= 16'h0176;    16'd31995: out <= 16'hFE15;
    16'd31996: out <= 16'hFAAE;    16'd31997: out <= 16'hFF00;    16'd31998: out <= 16'h0409;    16'd31999: out <= 16'hFD91;
    16'd32000: out <= 16'hFAAC;    16'd32001: out <= 16'hFE93;    16'd32002: out <= 16'h06D9;    16'd32003: out <= 16'hFF07;
    16'd32004: out <= 16'hFD2D;    16'd32005: out <= 16'hFF85;    16'd32006: out <= 16'hFD4D;    16'd32007: out <= 16'h0361;
    16'd32008: out <= 16'h0086;    16'd32009: out <= 16'hFE52;    16'd32010: out <= 16'h019D;    16'd32011: out <= 16'h0122;
    16'd32012: out <= 16'h0874;    16'd32013: out <= 16'hFC0A;    16'd32014: out <= 16'h0010;    16'd32015: out <= 16'hFE2E;
    16'd32016: out <= 16'h01C0;    16'd32017: out <= 16'h0730;    16'd32018: out <= 16'hFE9E;    16'd32019: out <= 16'hFA71;
    16'd32020: out <= 16'hFDA1;    16'd32021: out <= 16'h0255;    16'd32022: out <= 16'h01F6;    16'd32023: out <= 16'h0130;
    16'd32024: out <= 16'h0112;    16'd32025: out <= 16'h041E;    16'd32026: out <= 16'h0285;    16'd32027: out <= 16'hFEC4;
    16'd32028: out <= 16'hFC2B;    16'd32029: out <= 16'h03DF;    16'd32030: out <= 16'hFDF2;    16'd32031: out <= 16'h0734;
    16'd32032: out <= 16'h0263;    16'd32033: out <= 16'h0883;    16'd32034: out <= 16'hFDC2;    16'd32035: out <= 16'h0299;
    16'd32036: out <= 16'h056F;    16'd32037: out <= 16'h010D;    16'd32038: out <= 16'h02FF;    16'd32039: out <= 16'h0248;
    16'd32040: out <= 16'h0445;    16'd32041: out <= 16'h05B4;    16'd32042: out <= 16'h03FE;    16'd32043: out <= 16'h045F;
    16'd32044: out <= 16'h003A;    16'd32045: out <= 16'h0974;    16'd32046: out <= 16'h0E0F;    16'd32047: out <= 16'h049B;
    16'd32048: out <= 16'hF916;    16'd32049: out <= 16'h023A;    16'd32050: out <= 16'h043B;    16'd32051: out <= 16'h0551;
    16'd32052: out <= 16'h0023;    16'd32053: out <= 16'hFF5E;    16'd32054: out <= 16'h0571;    16'd32055: out <= 16'h02FF;
    16'd32056: out <= 16'h050A;    16'd32057: out <= 16'h04A9;    16'd32058: out <= 16'h0825;    16'd32059: out <= 16'h0023;
    16'd32060: out <= 16'h066E;    16'd32061: out <= 16'h04F0;    16'd32062: out <= 16'h046F;    16'd32063: out <= 16'h0103;
    16'd32064: out <= 16'h02A9;    16'd32065: out <= 16'h0731;    16'd32066: out <= 16'h069D;    16'd32067: out <= 16'h06E8;
    16'd32068: out <= 16'h04B0;    16'd32069: out <= 16'h0532;    16'd32070: out <= 16'h0104;    16'd32071: out <= 16'h0526;
    16'd32072: out <= 16'h00A1;    16'd32073: out <= 16'hFE32;    16'd32074: out <= 16'h000B;    16'd32075: out <= 16'h044E;
    16'd32076: out <= 16'h0355;    16'd32077: out <= 16'h04D4;    16'd32078: out <= 16'h055C;    16'd32079: out <= 16'h07AC;
    16'd32080: out <= 16'h01EB;    16'd32081: out <= 16'h0464;    16'd32082: out <= 16'h04F1;    16'd32083: out <= 16'h06D0;
    16'd32084: out <= 16'h01C0;    16'd32085: out <= 16'h00D2;    16'd32086: out <= 16'h07E6;    16'd32087: out <= 16'h0095;
    16'd32088: out <= 16'h0684;    16'd32089: out <= 16'h03A5;    16'd32090: out <= 16'h027F;    16'd32091: out <= 16'h0AF2;
    16'd32092: out <= 16'h025D;    16'd32093: out <= 16'h0298;    16'd32094: out <= 16'hF8B9;    16'd32095: out <= 16'h077B;
    16'd32096: out <= 16'hFFC0;    16'd32097: out <= 16'h07B9;    16'd32098: out <= 16'h0201;    16'd32099: out <= 16'hFCF2;
    16'd32100: out <= 16'h0290;    16'd32101: out <= 16'h058A;    16'd32102: out <= 16'hFFE9;    16'd32103: out <= 16'hFF88;
    16'd32104: out <= 16'hFFA9;    16'd32105: out <= 16'h031F;    16'd32106: out <= 16'h05DA;    16'd32107: out <= 16'h050F;
    16'd32108: out <= 16'h044D;    16'd32109: out <= 16'hFFB7;    16'd32110: out <= 16'h074E;    16'd32111: out <= 16'h097B;
    16'd32112: out <= 16'hFB66;    16'd32113: out <= 16'h01D2;    16'd32114: out <= 16'hFE24;    16'd32115: out <= 16'h0C2F;
    16'd32116: out <= 16'h08B2;    16'd32117: out <= 16'h07E7;    16'd32118: out <= 16'h07FC;    16'd32119: out <= 16'h076F;
    16'd32120: out <= 16'h076F;    16'd32121: out <= 16'h03ED;    16'd32122: out <= 16'h06AD;    16'd32123: out <= 16'h0060;
    16'd32124: out <= 16'h0810;    16'd32125: out <= 16'h06F1;    16'd32126: out <= 16'h058D;    16'd32127: out <= 16'h0854;
    16'd32128: out <= 16'h050C;    16'd32129: out <= 16'h0996;    16'd32130: out <= 16'h032C;    16'd32131: out <= 16'h02DB;
    16'd32132: out <= 16'hFFCD;    16'd32133: out <= 16'h01EE;    16'd32134: out <= 16'h0404;    16'd32135: out <= 16'h098A;
    16'd32136: out <= 16'h0853;    16'd32137: out <= 16'hFCE2;    16'd32138: out <= 16'hFBD4;    16'd32139: out <= 16'h0212;
    16'd32140: out <= 16'h0663;    16'd32141: out <= 16'h0614;    16'd32142: out <= 16'h0059;    16'd32143: out <= 16'h0506;
    16'd32144: out <= 16'h04A8;    16'd32145: out <= 16'h04D1;    16'd32146: out <= 16'hFF51;    16'd32147: out <= 16'h077B;
    16'd32148: out <= 16'h0BC6;    16'd32149: out <= 16'hFF0F;    16'd32150: out <= 16'h01E1;    16'd32151: out <= 16'hFF44;
    16'd32152: out <= 16'h03B5;    16'd32153: out <= 16'h0357;    16'd32154: out <= 16'h04CB;    16'd32155: out <= 16'h01D8;
    16'd32156: out <= 16'h0775;    16'd32157: out <= 16'h02A9;    16'd32158: out <= 16'h055F;    16'd32159: out <= 16'h03AF;
    16'd32160: out <= 16'h0394;    16'd32161: out <= 16'h00AE;    16'd32162: out <= 16'h08B9;    16'd32163: out <= 16'h0327;
    16'd32164: out <= 16'h0492;    16'd32165: out <= 16'h0408;    16'd32166: out <= 16'h0837;    16'd32167: out <= 16'h02F0;
    16'd32168: out <= 16'h01B0;    16'd32169: out <= 16'h0373;    16'd32170: out <= 16'h0830;    16'd32171: out <= 16'h059B;
    16'd32172: out <= 16'hFF66;    16'd32173: out <= 16'h0480;    16'd32174: out <= 16'h007D;    16'd32175: out <= 16'h062A;
    16'd32176: out <= 16'h04D2;    16'd32177: out <= 16'h02C3;    16'd32178: out <= 16'h0526;    16'd32179: out <= 16'h05CE;
    16'd32180: out <= 16'h07B9;    16'd32181: out <= 16'h0358;    16'd32182: out <= 16'h063F;    16'd32183: out <= 16'h0901;
    16'd32184: out <= 16'h077F;    16'd32185: out <= 16'h0080;    16'd32186: out <= 16'h03E6;    16'd32187: out <= 16'h02F7;
    16'd32188: out <= 16'h0A82;    16'd32189: out <= 16'hFD04;    16'd32190: out <= 16'h031C;    16'd32191: out <= 16'h033A;
    16'd32192: out <= 16'hFF04;    16'd32193: out <= 16'h0695;    16'd32194: out <= 16'h0E9C;    16'd32195: out <= 16'h016B;
    16'd32196: out <= 16'h0789;    16'd32197: out <= 16'hF8E9;    16'd32198: out <= 16'h091E;    16'd32199: out <= 16'hFFF4;
    16'd32200: out <= 16'h02CB;    16'd32201: out <= 16'h0F28;    16'd32202: out <= 16'h0389;    16'd32203: out <= 16'h03D8;
    16'd32204: out <= 16'h0F97;    16'd32205: out <= 16'h0776;    16'd32206: out <= 16'h0070;    16'd32207: out <= 16'h0023;
    16'd32208: out <= 16'h02EE;    16'd32209: out <= 16'h09FB;    16'd32210: out <= 16'h0B0F;    16'd32211: out <= 16'h0931;
    16'd32212: out <= 16'h058C;    16'd32213: out <= 16'h0D80;    16'd32214: out <= 16'h093C;    16'd32215: out <= 16'h0764;
    16'd32216: out <= 16'h08C5;    16'd32217: out <= 16'hFF87;    16'd32218: out <= 16'h027F;    16'd32219: out <= 16'h0570;
    16'd32220: out <= 16'hF9C5;    16'd32221: out <= 16'h0176;    16'd32222: out <= 16'h0379;    16'd32223: out <= 16'h0107;
    16'd32224: out <= 16'h0610;    16'd32225: out <= 16'hFFE0;    16'd32226: out <= 16'h032B;    16'd32227: out <= 16'h00DA;
    16'd32228: out <= 16'h084B;    16'd32229: out <= 16'h04DC;    16'd32230: out <= 16'hFCBF;    16'd32231: out <= 16'h018C;
    16'd32232: out <= 16'h05BF;    16'd32233: out <= 16'h0626;    16'd32234: out <= 16'hFAA6;    16'd32235: out <= 16'hFD3B;
    16'd32236: out <= 16'h0699;    16'd32237: out <= 16'h061B;    16'd32238: out <= 16'h03EC;    16'd32239: out <= 16'hFF1D;
    16'd32240: out <= 16'h0551;    16'd32241: out <= 16'hFC33;    16'd32242: out <= 16'h0706;    16'd32243: out <= 16'h014F;
    16'd32244: out <= 16'hFFB8;    16'd32245: out <= 16'hFF67;    16'd32246: out <= 16'h00EE;    16'd32247: out <= 16'hFBDE;
    16'd32248: out <= 16'hFDF8;    16'd32249: out <= 16'h0398;    16'd32250: out <= 16'hFDC1;    16'd32251: out <= 16'h0027;
    16'd32252: out <= 16'h0235;    16'd32253: out <= 16'hFB51;    16'd32254: out <= 16'h023A;    16'd32255: out <= 16'hFDF2;
    16'd32256: out <= 16'hFFAC;    16'd32257: out <= 16'h034C;    16'd32258: out <= 16'h0386;    16'd32259: out <= 16'h0495;
    16'd32260: out <= 16'h0420;    16'd32261: out <= 16'h027A;    16'd32262: out <= 16'hFADA;    16'd32263: out <= 16'hFD7B;
    16'd32264: out <= 16'hFC58;    16'd32265: out <= 16'hFEC9;    16'd32266: out <= 16'h0432;    16'd32267: out <= 16'hFEB3;
    16'd32268: out <= 16'h010A;    16'd32269: out <= 16'h0201;    16'd32270: out <= 16'hFE7A;    16'd32271: out <= 16'h01F9;
    16'd32272: out <= 16'hFF3D;    16'd32273: out <= 16'hFC14;    16'd32274: out <= 16'h004E;    16'd32275: out <= 16'h028E;
    16'd32276: out <= 16'h0101;    16'd32277: out <= 16'hFDEC;    16'd32278: out <= 16'hF790;    16'd32279: out <= 16'h0166;
    16'd32280: out <= 16'h00AA;    16'd32281: out <= 16'h0904;    16'd32282: out <= 16'h0709;    16'd32283: out <= 16'h0185;
    16'd32284: out <= 16'h041F;    16'd32285: out <= 16'hFFFA;    16'd32286: out <= 16'h0509;    16'd32287: out <= 16'h07A9;
    16'd32288: out <= 16'h0586;    16'd32289: out <= 16'h0321;    16'd32290: out <= 16'h01AE;    16'd32291: out <= 16'h01D7;
    16'd32292: out <= 16'h0529;    16'd32293: out <= 16'h035F;    16'd32294: out <= 16'h0553;    16'd32295: out <= 16'h061E;
    16'd32296: out <= 16'h07F7;    16'd32297: out <= 16'h0AA1;    16'd32298: out <= 16'h056D;    16'd32299: out <= 16'h0058;
    16'd32300: out <= 16'hFF76;    16'd32301: out <= 16'h0856;    16'd32302: out <= 16'h057F;    16'd32303: out <= 16'h0779;
    16'd32304: out <= 16'h044A;    16'd32305: out <= 16'h07FD;    16'd32306: out <= 16'h0196;    16'd32307: out <= 16'h0690;
    16'd32308: out <= 16'hFFD5;    16'd32309: out <= 16'hFCEC;    16'd32310: out <= 16'h097D;    16'd32311: out <= 16'h0624;
    16'd32312: out <= 16'h0760;    16'd32313: out <= 16'h063A;    16'd32314: out <= 16'h012C;    16'd32315: out <= 16'h0225;
    16'd32316: out <= 16'h0468;    16'd32317: out <= 16'h0216;    16'd32318: out <= 16'hFD50;    16'd32319: out <= 16'h020D;
    16'd32320: out <= 16'h00C1;    16'd32321: out <= 16'h01AA;    16'd32322: out <= 16'h068D;    16'd32323: out <= 16'h022D;
    16'd32324: out <= 16'hFF04;    16'd32325: out <= 16'h04D6;    16'd32326: out <= 16'h0A35;    16'd32327: out <= 16'h0556;
    16'd32328: out <= 16'h0A7B;    16'd32329: out <= 16'h05BE;    16'd32330: out <= 16'h050B;    16'd32331: out <= 16'h07D1;
    16'd32332: out <= 16'h022A;    16'd32333: out <= 16'h0901;    16'd32334: out <= 16'h00DB;    16'd32335: out <= 16'h1052;
    16'd32336: out <= 16'h0477;    16'd32337: out <= 16'h0585;    16'd32338: out <= 16'h040E;    16'd32339: out <= 16'hFB4C;
    16'd32340: out <= 16'h00BB;    16'd32341: out <= 16'h077D;    16'd32342: out <= 16'h0116;    16'd32343: out <= 16'hFE1E;
    16'd32344: out <= 16'h03CA;    16'd32345: out <= 16'h0649;    16'd32346: out <= 16'h00AF;    16'd32347: out <= 16'h0657;
    16'd32348: out <= 16'h03CE;    16'd32349: out <= 16'hFFDB;    16'd32350: out <= 16'h0367;    16'd32351: out <= 16'h0879;
    16'd32352: out <= 16'h0730;    16'd32353: out <= 16'hFEDB;    16'd32354: out <= 16'h04F9;    16'd32355: out <= 16'h0753;
    16'd32356: out <= 16'h011B;    16'd32357: out <= 16'h071D;    16'd32358: out <= 16'hFF76;    16'd32359: out <= 16'h0B34;
    16'd32360: out <= 16'h06BB;    16'd32361: out <= 16'h0495;    16'd32362: out <= 16'h006A;    16'd32363: out <= 16'h04C5;
    16'd32364: out <= 16'h0342;    16'd32365: out <= 16'h03DE;    16'd32366: out <= 16'h09F6;    16'd32367: out <= 16'hFEE8;
    16'd32368: out <= 16'h0800;    16'd32369: out <= 16'h01F2;    16'd32370: out <= 16'h0386;    16'd32371: out <= 16'h0625;
    16'd32372: out <= 16'h00C0;    16'd32373: out <= 16'hFEF3;    16'd32374: out <= 16'h0B73;    16'd32375: out <= 16'h03FD;
    16'd32376: out <= 16'h0BD8;    16'd32377: out <= 16'h03EF;    16'd32378: out <= 16'hFFF1;    16'd32379: out <= 16'h0118;
    16'd32380: out <= 16'hFD87;    16'd32381: out <= 16'h0390;    16'd32382: out <= 16'hFE3A;    16'd32383: out <= 16'h08EC;
    16'd32384: out <= 16'h0920;    16'd32385: out <= 16'h03EF;    16'd32386: out <= 16'h03C4;    16'd32387: out <= 16'h08D1;
    16'd32388: out <= 16'h0A78;    16'd32389: out <= 16'h020A;    16'd32390: out <= 16'h0211;    16'd32391: out <= 16'h0958;
    16'd32392: out <= 16'h0712;    16'd32393: out <= 16'h038A;    16'd32394: out <= 16'h033F;    16'd32395: out <= 16'h000C;
    16'd32396: out <= 16'hFE5C;    16'd32397: out <= 16'h09F9;    16'd32398: out <= 16'hFF92;    16'd32399: out <= 16'h02FA;
    16'd32400: out <= 16'hFC9E;    16'd32401: out <= 16'h0776;    16'd32402: out <= 16'h024B;    16'd32403: out <= 16'hFABD;
    16'd32404: out <= 16'h0443;    16'd32405: out <= 16'h024E;    16'd32406: out <= 16'h045D;    16'd32407: out <= 16'h05BB;
    16'd32408: out <= 16'h047C;    16'd32409: out <= 16'hFD5E;    16'd32410: out <= 16'hFCEA;    16'd32411: out <= 16'hFB3B;
    16'd32412: out <= 16'h07D0;    16'd32413: out <= 16'hFF36;    16'd32414: out <= 16'hFD0A;    16'd32415: out <= 16'h0116;
    16'd32416: out <= 16'h01FC;    16'd32417: out <= 16'h01A2;    16'd32418: out <= 16'hFDBB;    16'd32419: out <= 16'h01A2;
    16'd32420: out <= 16'h005C;    16'd32421: out <= 16'h017F;    16'd32422: out <= 16'h0673;    16'd32423: out <= 16'h048C;
    16'd32424: out <= 16'h0443;    16'd32425: out <= 16'h00C9;    16'd32426: out <= 16'hFAD6;    16'd32427: out <= 16'h0CC2;
    16'd32428: out <= 16'h042D;    16'd32429: out <= 16'h054E;    16'd32430: out <= 16'h08C5;    16'd32431: out <= 16'h02C8;
    16'd32432: out <= 16'h03EB;    16'd32433: out <= 16'h0382;    16'd32434: out <= 16'h018E;    16'd32435: out <= 16'h00ED;
    16'd32436: out <= 16'h019A;    16'd32437: out <= 16'h0ED5;    16'd32438: out <= 16'h0617;    16'd32439: out <= 16'hFEC9;
    16'd32440: out <= 16'h05B6;    16'd32441: out <= 16'hFBB0;    16'd32442: out <= 16'hFFCA;    16'd32443: out <= 16'h0769;
    16'd32444: out <= 16'h0872;    16'd32445: out <= 16'h08BF;    16'd32446: out <= 16'h01DB;    16'd32447: out <= 16'h0005;
    16'd32448: out <= 16'h028F;    16'd32449: out <= 16'h08DF;    16'd32450: out <= 16'h04E8;    16'd32451: out <= 16'h04DF;
    16'd32452: out <= 16'h04F2;    16'd32453: out <= 16'h05A6;    16'd32454: out <= 16'h0830;    16'd32455: out <= 16'h02F0;
    16'd32456: out <= 16'h01ED;    16'd32457: out <= 16'h0B32;    16'd32458: out <= 16'h0377;    16'd32459: out <= 16'h05F2;
    16'd32460: out <= 16'h05F5;    16'd32461: out <= 16'hFFC3;    16'd32462: out <= 16'hFEBC;    16'd32463: out <= 16'h015F;
    16'd32464: out <= 16'h029B;    16'd32465: out <= 16'h05CB;    16'd32466: out <= 16'hFEF7;    16'd32467: out <= 16'h008C;
    16'd32468: out <= 16'h0326;    16'd32469: out <= 16'h0066;    16'd32470: out <= 16'h0290;    16'd32471: out <= 16'hF99F;
    16'd32472: out <= 16'h0514;    16'd32473: out <= 16'hFD20;    16'd32474: out <= 16'h040A;    16'd32475: out <= 16'h000F;
    16'd32476: out <= 16'h0AE2;    16'd32477: out <= 16'h025B;    16'd32478: out <= 16'h024C;    16'd32479: out <= 16'hFF11;
    16'd32480: out <= 16'h0643;    16'd32481: out <= 16'h0209;    16'd32482: out <= 16'h03B9;    16'd32483: out <= 16'h0217;
    16'd32484: out <= 16'h0C6F;    16'd32485: out <= 16'h00E8;    16'd32486: out <= 16'h05FC;    16'd32487: out <= 16'h02F4;
    16'd32488: out <= 16'h0136;    16'd32489: out <= 16'hFDCD;    16'd32490: out <= 16'h025B;    16'd32491: out <= 16'h045A;
    16'd32492: out <= 16'hFC73;    16'd32493: out <= 16'h049B;    16'd32494: out <= 16'hFB69;    16'd32495: out <= 16'hFBDB;
    16'd32496: out <= 16'h0435;    16'd32497: out <= 16'h06BC;    16'd32498: out <= 16'h0037;    16'd32499: out <= 16'h02F3;
    16'd32500: out <= 16'hFDE4;    16'd32501: out <= 16'h014B;    16'd32502: out <= 16'hFCB6;    16'd32503: out <= 16'hF6AC;
    16'd32504: out <= 16'h0197;    16'd32505: out <= 16'hFFA4;    16'd32506: out <= 16'hFD4B;    16'd32507: out <= 16'hFE98;
    16'd32508: out <= 16'hFFB9;    16'd32509: out <= 16'h031F;    16'd32510: out <= 16'h035E;    16'd32511: out <= 16'hFBE8;
    16'd32512: out <= 16'h06DC;    16'd32513: out <= 16'h0529;    16'd32514: out <= 16'hFF27;    16'd32515: out <= 16'hFD52;
    16'd32516: out <= 16'hFD7C;    16'd32517: out <= 16'h05F5;    16'd32518: out <= 16'hFF9B;    16'd32519: out <= 16'h01E7;
    16'd32520: out <= 16'hFD00;    16'd32521: out <= 16'hFF12;    16'd32522: out <= 16'h0394;    16'd32523: out <= 16'h0222;
    16'd32524: out <= 16'h0163;    16'd32525: out <= 16'h00BF;    16'd32526: out <= 16'h06EA;    16'd32527: out <= 16'hFE4C;
    16'd32528: out <= 16'hFCC1;    16'd32529: out <= 16'hFE24;    16'd32530: out <= 16'hFA5E;    16'd32531: out <= 16'h0424;
    16'd32532: out <= 16'h05F6;    16'd32533: out <= 16'hFAB6;    16'd32534: out <= 16'h02DC;    16'd32535: out <= 16'h07AC;
    16'd32536: out <= 16'hFEE5;    16'd32537: out <= 16'h05DB;    16'd32538: out <= 16'hFF46;    16'd32539: out <= 16'h0568;
    16'd32540: out <= 16'hFB04;    16'd32541: out <= 16'h0318;    16'd32542: out <= 16'h07EE;    16'd32543: out <= 16'h02FA;
    16'd32544: out <= 16'h097C;    16'd32545: out <= 16'h00BB;    16'd32546: out <= 16'h082E;    16'd32547: out <= 16'h06C2;
    16'd32548: out <= 16'h03C9;    16'd32549: out <= 16'h090F;    16'd32550: out <= 16'h021A;    16'd32551: out <= 16'h0479;
    16'd32552: out <= 16'h00C1;    16'd32553: out <= 16'h011F;    16'd32554: out <= 16'h0751;    16'd32555: out <= 16'h04DE;
    16'd32556: out <= 16'h036B;    16'd32557: out <= 16'h0674;    16'd32558: out <= 16'h0292;    16'd32559: out <= 16'h03FE;
    16'd32560: out <= 16'h05BA;    16'd32561: out <= 16'h02D4;    16'd32562: out <= 16'h031B;    16'd32563: out <= 16'h03B6;
    16'd32564: out <= 16'h05B2;    16'd32565: out <= 16'h060C;    16'd32566: out <= 16'h02AD;    16'd32567: out <= 16'hFB21;
    16'd32568: out <= 16'h01CB;    16'd32569: out <= 16'h072B;    16'd32570: out <= 16'h0345;    16'd32571: out <= 16'h097B;
    16'd32572: out <= 16'h09A8;    16'd32573: out <= 16'h0B82;    16'd32574: out <= 16'h0B8A;    16'd32575: out <= 16'h0D8E;
    16'd32576: out <= 16'h029E;    16'd32577: out <= 16'h0521;    16'd32578: out <= 16'h0444;    16'd32579: out <= 16'h00F0;
    16'd32580: out <= 16'h0899;    16'd32581: out <= 16'h0AB8;    16'd32582: out <= 16'h03C8;    16'd32583: out <= 16'hFDD1;
    16'd32584: out <= 16'h03E0;    16'd32585: out <= 16'h03F9;    16'd32586: out <= 16'h095C;    16'd32587: out <= 16'h0688;
    16'd32588: out <= 16'h043F;    16'd32589: out <= 16'h00AC;    16'd32590: out <= 16'h00E2;    16'd32591: out <= 16'h0060;
    16'd32592: out <= 16'h0736;    16'd32593: out <= 16'h0469;    16'd32594: out <= 16'h0606;    16'd32595: out <= 16'hFFE9;
    16'd32596: out <= 16'h02A1;    16'd32597: out <= 16'h0644;    16'd32598: out <= 16'h0485;    16'd32599: out <= 16'h0768;
    16'd32600: out <= 16'h0630;    16'd32601: out <= 16'hFE98;    16'd32602: out <= 16'hFC7D;    16'd32603: out <= 16'h0188;
    16'd32604: out <= 16'h01FE;    16'd32605: out <= 16'h0A77;    16'd32606: out <= 16'h0580;    16'd32607: out <= 16'h06E1;
    16'd32608: out <= 16'h00DB;    16'd32609: out <= 16'h081D;    16'd32610: out <= 16'hFC61;    16'd32611: out <= 16'h0A92;
    16'd32612: out <= 16'h07DA;    16'd32613: out <= 16'h02F2;    16'd32614: out <= 16'h061E;    16'd32615: out <= 16'h0E91;
    16'd32616: out <= 16'h004B;    16'd32617: out <= 16'h0786;    16'd32618: out <= 16'h08CD;    16'd32619: out <= 16'h03D2;
    16'd32620: out <= 16'h06FE;    16'd32621: out <= 16'h0473;    16'd32622: out <= 16'h0294;    16'd32623: out <= 16'h0D1D;
    16'd32624: out <= 16'h0641;    16'd32625: out <= 16'h05DA;    16'd32626: out <= 16'h0527;    16'd32627: out <= 16'h0C6E;
    16'd32628: out <= 16'h05E7;    16'd32629: out <= 16'h12D8;    16'd32630: out <= 16'h002E;    16'd32631: out <= 16'hFD67;
    16'd32632: out <= 16'hFF61;    16'd32633: out <= 16'h0A8E;    16'd32634: out <= 16'h09F2;    16'd32635: out <= 16'h088E;
    16'd32636: out <= 16'h0642;    16'd32637: out <= 16'h040C;    16'd32638: out <= 16'h0589;    16'd32639: out <= 16'h0938;
    16'd32640: out <= 16'h0B53;    16'd32641: out <= 16'hFFE9;    16'd32642: out <= 16'h071B;    16'd32643: out <= 16'h00EB;
    16'd32644: out <= 16'h0578;    16'd32645: out <= 16'h09BE;    16'd32646: out <= 16'h05DE;    16'd32647: out <= 16'h09B1;
    16'd32648: out <= 16'h00BD;    16'd32649: out <= 16'h0151;    16'd32650: out <= 16'h06EC;    16'd32651: out <= 16'hFF82;
    16'd32652: out <= 16'h03F4;    16'd32653: out <= 16'h0578;    16'd32654: out <= 16'h03E8;    16'd32655: out <= 16'hFE8F;
    16'd32656: out <= 16'hFE8E;    16'd32657: out <= 16'h0212;    16'd32658: out <= 16'h06B0;    16'd32659: out <= 16'h068B;
    16'd32660: out <= 16'h01F1;    16'd32661: out <= 16'h0877;    16'd32662: out <= 16'h03F2;    16'd32663: out <= 16'hFEEB;
    16'd32664: out <= 16'h0A8A;    16'd32665: out <= 16'hFFD6;    16'd32666: out <= 16'h08CD;    16'd32667: out <= 16'h0184;
    16'd32668: out <= 16'h08CA;    16'd32669: out <= 16'h0928;    16'd32670: out <= 16'h042A;    16'd32671: out <= 16'hFD8C;
    16'd32672: out <= 16'h048F;    16'd32673: out <= 16'h05E3;    16'd32674: out <= 16'h00FC;    16'd32675: out <= 16'hFF8F;
    16'd32676: out <= 16'h0288;    16'd32677: out <= 16'h0390;    16'd32678: out <= 16'h082E;    16'd32679: out <= 16'h0B0D;
    16'd32680: out <= 16'h0358;    16'd32681: out <= 16'h05A4;    16'd32682: out <= 16'hFF0F;    16'd32683: out <= 16'hFEE9;
    16'd32684: out <= 16'h058B;    16'd32685: out <= 16'h022A;    16'd32686: out <= 16'h01D8;    16'd32687: out <= 16'h02D2;
    16'd32688: out <= 16'h0226;    16'd32689: out <= 16'h093F;    16'd32690: out <= 16'h12CA;    16'd32691: out <= 16'h0612;
    16'd32692: out <= 16'h0092;    16'd32693: out <= 16'h0203;    16'd32694: out <= 16'h049F;    16'd32695: out <= 16'h078E;
    16'd32696: out <= 16'h0373;    16'd32697: out <= 16'hFD5C;    16'd32698: out <= 16'hFE28;    16'd32699: out <= 16'h08E3;
    16'd32700: out <= 16'h056D;    16'd32701: out <= 16'hFD33;    16'd32702: out <= 16'h056C;    16'd32703: out <= 16'h06EE;
    16'd32704: out <= 16'hFE02;    16'd32705: out <= 16'h04C5;    16'd32706: out <= 16'h0E9C;    16'd32707: out <= 16'h064C;
    16'd32708: out <= 16'h0AE1;    16'd32709: out <= 16'h07B2;    16'd32710: out <= 16'h0173;    16'd32711: out <= 16'h02E6;
    16'd32712: out <= 16'hFF8D;    16'd32713: out <= 16'h07A7;    16'd32714: out <= 16'h0B68;    16'd32715: out <= 16'h0DB9;
    16'd32716: out <= 16'h0739;    16'd32717: out <= 16'h038F;    16'd32718: out <= 16'hFDF6;    16'd32719: out <= 16'h07E8;
    16'd32720: out <= 16'h0475;    16'd32721: out <= 16'h0541;    16'd32722: out <= 16'h0313;    16'd32723: out <= 16'h03B7;
    16'd32724: out <= 16'h06C3;    16'd32725: out <= 16'h0313;    16'd32726: out <= 16'hFE2A;    16'd32727: out <= 16'h05D9;
    16'd32728: out <= 16'h0252;    16'd32729: out <= 16'h01BC;    16'd32730: out <= 16'hFEAE;    16'd32731: out <= 16'hFCA2;
    16'd32732: out <= 16'h0556;    16'd32733: out <= 16'h0285;    16'd32734: out <= 16'h036F;    16'd32735: out <= 16'hFE00;
    16'd32736: out <= 16'h031D;    16'd32737: out <= 16'h08C9;    16'd32738: out <= 16'h0575;    16'd32739: out <= 16'h00BC;
    16'd32740: out <= 16'h0B19;    16'd32741: out <= 16'h049F;    16'd32742: out <= 16'hFB28;    16'd32743: out <= 16'h007F;
    16'd32744: out <= 16'hFF4A;    16'd32745: out <= 16'h0745;    16'd32746: out <= 16'hFCA1;    16'd32747: out <= 16'hFBF8;
    16'd32748: out <= 16'hFE7A;    16'd32749: out <= 16'hFDA6;    16'd32750: out <= 16'hFEE6;    16'd32751: out <= 16'hFF69;
    16'd32752: out <= 16'hFEB9;    16'd32753: out <= 16'h03C5;    16'd32754: out <= 16'hFE03;    16'd32755: out <= 16'h0017;
    16'd32756: out <= 16'hFE06;    16'd32757: out <= 16'h0799;    16'd32758: out <= 16'hFEC6;    16'd32759: out <= 16'hFD17;
    16'd32760: out <= 16'h0483;    16'd32761: out <= 16'h0340;    16'd32762: out <= 16'hF6FB;    16'd32763: out <= 16'h07BA;
    16'd32764: out <= 16'hFB2D;    16'd32765: out <= 16'hFCC5;    16'd32766: out <= 16'h0BB7;    16'd32767: out <= 16'h0015;
    16'd32768: out <= 16'h0150;    16'd32769: out <= 16'h04E8;    16'd32770: out <= 16'h01FB;    16'd32771: out <= 16'hFFE6;
    16'd32772: out <= 16'h0472;    16'd32773: out <= 16'hFD70;    16'd32774: out <= 16'h040F;    16'd32775: out <= 16'hFE98;
    16'd32776: out <= 16'hFDE7;    16'd32777: out <= 16'h0110;    16'd32778: out <= 16'h0117;    16'd32779: out <= 16'hFDA9;
    16'd32780: out <= 16'hFE14;    16'd32781: out <= 16'h0168;    16'd32782: out <= 16'h02D4;    16'd32783: out <= 16'hFABA;
    16'd32784: out <= 16'h0112;    16'd32785: out <= 16'h0041;    16'd32786: out <= 16'hFB7A;    16'd32787: out <= 16'h0372;
    16'd32788: out <= 16'h0570;    16'd32789: out <= 16'hFD75;    16'd32790: out <= 16'hFD6E;    16'd32791: out <= 16'h0067;
    16'd32792: out <= 16'h0619;    16'd32793: out <= 16'h0BEC;    16'd32794: out <= 16'h01D7;    16'd32795: out <= 16'hFFA1;
    16'd32796: out <= 16'hFE03;    16'd32797: out <= 16'h05CC;    16'd32798: out <= 16'h0363;    16'd32799: out <= 16'h081F;
    16'd32800: out <= 16'hFE4C;    16'd32801: out <= 16'h0936;    16'd32802: out <= 16'h06DF;    16'd32803: out <= 16'h01AF;
    16'd32804: out <= 16'h030D;    16'd32805: out <= 16'h04EB;    16'd32806: out <= 16'h05EC;    16'd32807: out <= 16'h0162;
    16'd32808: out <= 16'h0319;    16'd32809: out <= 16'h0811;    16'd32810: out <= 16'h00E1;    16'd32811: out <= 16'h05AD;
    16'd32812: out <= 16'h021A;    16'd32813: out <= 16'h0587;    16'd32814: out <= 16'h0926;    16'd32815: out <= 16'h03AB;
    16'd32816: out <= 16'h0670;    16'd32817: out <= 16'h03F8;    16'd32818: out <= 16'h058E;    16'd32819: out <= 16'h01E0;
    16'd32820: out <= 16'h0801;    16'd32821: out <= 16'h037F;    16'd32822: out <= 16'h0640;    16'd32823: out <= 16'h0127;
    16'd32824: out <= 16'h07ED;    16'd32825: out <= 16'h0292;    16'd32826: out <= 16'h0482;    16'd32827: out <= 16'h0D80;
    16'd32828: out <= 16'hFDE1;    16'd32829: out <= 16'h0288;    16'd32830: out <= 16'h011A;    16'd32831: out <= 16'hFF2B;
    16'd32832: out <= 16'h046C;    16'd32833: out <= 16'h02FC;    16'd32834: out <= 16'h06B3;    16'd32835: out <= 16'h0536;
    16'd32836: out <= 16'hFED6;    16'd32837: out <= 16'h0004;    16'd32838: out <= 16'hFDB5;    16'd32839: out <= 16'hFFF5;
    16'd32840: out <= 16'h05B8;    16'd32841: out <= 16'h0258;    16'd32842: out <= 16'h08D3;    16'd32843: out <= 16'h07E6;
    16'd32844: out <= 16'hFCFA;    16'd32845: out <= 16'hFF58;    16'd32846: out <= 16'h0760;    16'd32847: out <= 16'h011A;
    16'd32848: out <= 16'h070B;    16'd32849: out <= 16'h02B8;    16'd32850: out <= 16'h0A9A;    16'd32851: out <= 16'h024C;
    16'd32852: out <= 16'hFF62;    16'd32853: out <= 16'h05FF;    16'd32854: out <= 16'h0B73;    16'd32855: out <= 16'h0965;
    16'd32856: out <= 16'h0299;    16'd32857: out <= 16'h0501;    16'd32858: out <= 16'h07AB;    16'd32859: out <= 16'h03E5;
    16'd32860: out <= 16'h0274;    16'd32861: out <= 16'hFCA7;    16'd32862: out <= 16'h0376;    16'd32863: out <= 16'hF493;
    16'd32864: out <= 16'h09DE;    16'd32865: out <= 16'h00FB;    16'd32866: out <= 16'h0B06;    16'd32867: out <= 16'h01EA;
    16'd32868: out <= 16'h0247;    16'd32869: out <= 16'h06E5;    16'd32870: out <= 16'h0600;    16'd32871: out <= 16'h0CB6;
    16'd32872: out <= 16'hF82B;    16'd32873: out <= 16'h02DE;    16'd32874: out <= 16'h033D;    16'd32875: out <= 16'h07E5;
    16'd32876: out <= 16'h05E8;    16'd32877: out <= 16'hF9F1;    16'd32878: out <= 16'h067A;    16'd32879: out <= 16'h06DB;
    16'd32880: out <= 16'hFF8A;    16'd32881: out <= 16'h061A;    16'd32882: out <= 16'h01FB;    16'd32883: out <= 16'h0138;
    16'd32884: out <= 16'h0491;    16'd32885: out <= 16'h0667;    16'd32886: out <= 16'h061C;    16'd32887: out <= 16'h07BC;
    16'd32888: out <= 16'h022C;    16'd32889: out <= 16'hFEF2;    16'd32890: out <= 16'h0917;    16'd32891: out <= 16'h0CBD;
    16'd32892: out <= 16'h045E;    16'd32893: out <= 16'hFE9C;    16'd32894: out <= 16'hFE0C;    16'd32895: out <= 16'h0570;
    16'd32896: out <= 16'hFE3E;    16'd32897: out <= 16'h02D8;    16'd32898: out <= 16'h0303;    16'd32899: out <= 16'h043A;
    16'd32900: out <= 16'h0516;    16'd32901: out <= 16'h0257;    16'd32902: out <= 16'h00C3;    16'd32903: out <= 16'h0495;
    16'd32904: out <= 16'h0586;    16'd32905: out <= 16'hFB49;    16'd32906: out <= 16'h0137;    16'd32907: out <= 16'h03F2;
    16'd32908: out <= 16'h052F;    16'd32909: out <= 16'h05F0;    16'd32910: out <= 16'h00EA;    16'd32911: out <= 16'h064D;
    16'd32912: out <= 16'h05CC;    16'd32913: out <= 16'h04C0;    16'd32914: out <= 16'h023E;    16'd32915: out <= 16'h034C;
    16'd32916: out <= 16'h0407;    16'd32917: out <= 16'h033C;    16'd32918: out <= 16'h01F5;    16'd32919: out <= 16'h0398;
    16'd32920: out <= 16'h0AF1;    16'd32921: out <= 16'h04E1;    16'd32922: out <= 16'hFBCF;    16'd32923: out <= 16'h092C;
    16'd32924: out <= 16'h0523;    16'd32925: out <= 16'h04F2;    16'd32926: out <= 16'h0877;    16'd32927: out <= 16'h0372;
    16'd32928: out <= 16'h0408;    16'd32929: out <= 16'h0248;    16'd32930: out <= 16'h0B16;    16'd32931: out <= 16'h017E;
    16'd32932: out <= 16'h0303;    16'd32933: out <= 16'h0A4C;    16'd32934: out <= 16'h01ED;    16'd32935: out <= 16'h0439;
    16'd32936: out <= 16'h0229;    16'd32937: out <= 16'hFE95;    16'd32938: out <= 16'h0112;    16'd32939: out <= 16'h01E8;
    16'd32940: out <= 16'h04A1;    16'd32941: out <= 16'hFC35;    16'd32942: out <= 16'h037A;    16'd32943: out <= 16'h03D1;
    16'd32944: out <= 16'h07DE;    16'd32945: out <= 16'h01D1;    16'd32946: out <= 16'h0169;    16'd32947: out <= 16'h0274;
    16'd32948: out <= 16'h097D;    16'd32949: out <= 16'h081C;    16'd32950: out <= 16'h056C;    16'd32951: out <= 16'h054D;
    16'd32952: out <= 16'h02F9;    16'd32953: out <= 16'h0B20;    16'd32954: out <= 16'h0181;    16'd32955: out <= 16'h0371;
    16'd32956: out <= 16'h07BE;    16'd32957: out <= 16'h06EC;    16'd32958: out <= 16'hFF36;    16'd32959: out <= 16'h0A2C;
    16'd32960: out <= 16'h0391;    16'd32961: out <= 16'h03BD;    16'd32962: out <= 16'h0031;    16'd32963: out <= 16'h0C9C;
    16'd32964: out <= 16'h0490;    16'd32965: out <= 16'h04C0;    16'd32966: out <= 16'h03A4;    16'd32967: out <= 16'h012F;
    16'd32968: out <= 16'h0465;    16'd32969: out <= 16'h0477;    16'd32970: out <= 16'h087C;    16'd32971: out <= 16'h072F;
    16'd32972: out <= 16'hFDB1;    16'd32973: out <= 16'h00DA;    16'd32974: out <= 16'h0893;    16'd32975: out <= 16'h0385;
    16'd32976: out <= 16'hFF07;    16'd32977: out <= 16'hFE12;    16'd32978: out <= 16'h0764;    16'd32979: out <= 16'hFD46;
    16'd32980: out <= 16'h0153;    16'd32981: out <= 16'h05C0;    16'd32982: out <= 16'hFB88;    16'd32983: out <= 16'hFF94;
    16'd32984: out <= 16'hFE31;    16'd32985: out <= 16'hFB8F;    16'd32986: out <= 16'hFCCC;    16'd32987: out <= 16'h00DF;
    16'd32988: out <= 16'h094F;    16'd32989: out <= 16'h0526;    16'd32990: out <= 16'hFFE5;    16'd32991: out <= 16'h09C3;
    16'd32992: out <= 16'h0A4B;    16'd32993: out <= 16'h07AA;    16'd32994: out <= 16'h05EA;    16'd32995: out <= 16'h0430;
    16'd32996: out <= 16'h09B6;    16'd32997: out <= 16'h0923;    16'd32998: out <= 16'h056D;    16'd32999: out <= 16'hFB5F;
    16'd33000: out <= 16'h02B8;    16'd33001: out <= 16'h0835;    16'd33002: out <= 16'h0575;    16'd33003: out <= 16'h0513;
    16'd33004: out <= 16'hFBEA;    16'd33005: out <= 16'hFDBE;    16'd33006: out <= 16'hFE4C;    16'd33007: out <= 16'hFE12;
    16'd33008: out <= 16'h0321;    16'd33009: out <= 16'hFF0B;    16'd33010: out <= 16'hF7C0;    16'd33011: out <= 16'h0001;
    16'd33012: out <= 16'h018E;    16'd33013: out <= 16'h00E9;    16'd33014: out <= 16'hFD69;    16'd33015: out <= 16'hFE92;
    16'd33016: out <= 16'hFD9B;    16'd33017: out <= 16'h04CC;    16'd33018: out <= 16'h0670;    16'd33019: out <= 16'hFEC4;
    16'd33020: out <= 16'h0102;    16'd33021: out <= 16'hFB2E;    16'd33022: out <= 16'h02FB;    16'd33023: out <= 16'hFCF4;
    16'd33024: out <= 16'hFDD5;    16'd33025: out <= 16'hFFE0;    16'd33026: out <= 16'hFEA5;    16'd33027: out <= 16'hF83C;
    16'd33028: out <= 16'hFDED;    16'd33029: out <= 16'h07AA;    16'd33030: out <= 16'hFE18;    16'd33031: out <= 16'hFD38;
    16'd33032: out <= 16'h00C4;    16'd33033: out <= 16'h040D;    16'd33034: out <= 16'hFC40;    16'd33035: out <= 16'hF700;
    16'd33036: out <= 16'hFEA9;    16'd33037: out <= 16'h0999;    16'd33038: out <= 16'hFF70;    16'd33039: out <= 16'hFBE3;
    16'd33040: out <= 16'h034C;    16'd33041: out <= 16'h01A6;    16'd33042: out <= 16'hFDB7;    16'd33043: out <= 16'hFDC8;
    16'd33044: out <= 16'hFFC0;    16'd33045: out <= 16'hFF7D;    16'd33046: out <= 16'h0B0F;    16'd33047: out <= 16'h08C3;
    16'd33048: out <= 16'h0728;    16'd33049: out <= 16'h06CD;    16'd33050: out <= 16'h0911;    16'd33051: out <= 16'hFECE;
    16'd33052: out <= 16'hFCBA;    16'd33053: out <= 16'h043A;    16'd33054: out <= 16'hFEE4;    16'd33055: out <= 16'h01DD;
    16'd33056: out <= 16'hFEF9;    16'd33057: out <= 16'h0028;    16'd33058: out <= 16'h03FC;    16'd33059: out <= 16'h05AB;
    16'd33060: out <= 16'h01DA;    16'd33061: out <= 16'h03AB;    16'd33062: out <= 16'h0796;    16'd33063: out <= 16'h0824;
    16'd33064: out <= 16'h01A3;    16'd33065: out <= 16'hFDE8;    16'd33066: out <= 16'h0142;    16'd33067: out <= 16'h044C;
    16'd33068: out <= 16'h0298;    16'd33069: out <= 16'h0966;    16'd33070: out <= 16'h07BB;    16'd33071: out <= 16'h07D9;
    16'd33072: out <= 16'h03BE;    16'd33073: out <= 16'h0AC0;    16'd33074: out <= 16'h017D;    16'd33075: out <= 16'h0606;
    16'd33076: out <= 16'h0293;    16'd33077: out <= 16'h06D4;    16'd33078: out <= 16'h000D;    16'd33079: out <= 16'h04CD;
    16'd33080: out <= 16'h0132;    16'd33081: out <= 16'h03D4;    16'd33082: out <= 16'hFCF7;    16'd33083: out <= 16'h01F2;
    16'd33084: out <= 16'h02A3;    16'd33085: out <= 16'h059B;    16'd33086: out <= 16'hFF40;    16'd33087: out <= 16'h06AC;
    16'd33088: out <= 16'hFE0F;    16'd33089: out <= 16'h090D;    16'd33090: out <= 16'hFC96;    16'd33091: out <= 16'h006A;
    16'd33092: out <= 16'hFF0C;    16'd33093: out <= 16'h02A0;    16'd33094: out <= 16'h02DC;    16'd33095: out <= 16'h0179;
    16'd33096: out <= 16'h0554;    16'd33097: out <= 16'hFDCF;    16'd33098: out <= 16'h05DD;    16'd33099: out <= 16'h0275;
    16'd33100: out <= 16'h0226;    16'd33101: out <= 16'h0AB6;    16'd33102: out <= 16'h00A8;    16'd33103: out <= 16'h024E;
    16'd33104: out <= 16'h04D2;    16'd33105: out <= 16'h0946;    16'd33106: out <= 16'h00FB;    16'd33107: out <= 16'h0904;
    16'd33108: out <= 16'h0497;    16'd33109: out <= 16'h046D;    16'd33110: out <= 16'h0484;    16'd33111: out <= 16'h01CF;
    16'd33112: out <= 16'h046F;    16'd33113: out <= 16'h03EE;    16'd33114: out <= 16'h03BB;    16'd33115: out <= 16'h0656;
    16'd33116: out <= 16'h0287;    16'd33117: out <= 16'h05A9;    16'd33118: out <= 16'hFD97;    16'd33119: out <= 16'h0B38;
    16'd33120: out <= 16'h019E;    16'd33121: out <= 16'h08C5;    16'd33122: out <= 16'h03BB;    16'd33123: out <= 16'hFFC4;
    16'd33124: out <= 16'h0522;    16'd33125: out <= 16'hFE44;    16'd33126: out <= 16'h0031;    16'd33127: out <= 16'h039C;
    16'd33128: out <= 16'hFB89;    16'd33129: out <= 16'h0E3C;    16'd33130: out <= 16'h0272;    16'd33131: out <= 16'h04A9;
    16'd33132: out <= 16'h07F6;    16'd33133: out <= 16'h0178;    16'd33134: out <= 16'h0A74;    16'd33135: out <= 16'h0B20;
    16'd33136: out <= 16'hFF00;    16'd33137: out <= 16'h06E7;    16'd33138: out <= 16'h0155;    16'd33139: out <= 16'h0621;
    16'd33140: out <= 16'h06AF;    16'd33141: out <= 16'h0077;    16'd33142: out <= 16'h0505;    16'd33143: out <= 16'h06F6;
    16'd33144: out <= 16'hFEAF;    16'd33145: out <= 16'hFD77;    16'd33146: out <= 16'h04AB;    16'd33147: out <= 16'h0130;
    16'd33148: out <= 16'h04D6;    16'd33149: out <= 16'h0825;    16'd33150: out <= 16'hFEB8;    16'd33151: out <= 16'h0384;
    16'd33152: out <= 16'h0636;    16'd33153: out <= 16'h0201;    16'd33154: out <= 16'h02B7;    16'd33155: out <= 16'hFC08;
    16'd33156: out <= 16'h0265;    16'd33157: out <= 16'h03D8;    16'd33158: out <= 16'h0AB4;    16'd33159: out <= 16'h01B4;
    16'd33160: out <= 16'h0258;    16'd33161: out <= 16'h0EB7;    16'd33162: out <= 16'h02FC;    16'd33163: out <= 16'h07EB;
    16'd33164: out <= 16'h0783;    16'd33165: out <= 16'hFEB4;    16'd33166: out <= 16'h02C7;    16'd33167: out <= 16'h006E;
    16'd33168: out <= 16'h00FA;    16'd33169: out <= 16'h06FE;    16'd33170: out <= 16'h083C;    16'd33171: out <= 16'h0BA6;
    16'd33172: out <= 16'hFED3;    16'd33173: out <= 16'h05D1;    16'd33174: out <= 16'hFECF;    16'd33175: out <= 16'h0555;
    16'd33176: out <= 16'h07B4;    16'd33177: out <= 16'h0593;    16'd33178: out <= 16'hF9BD;    16'd33179: out <= 16'h01F6;
    16'd33180: out <= 16'h01AF;    16'd33181: out <= 16'h0B35;    16'd33182: out <= 16'h053B;    16'd33183: out <= 16'h0358;
    16'd33184: out <= 16'h0565;    16'd33185: out <= 16'hFEFF;    16'd33186: out <= 16'hFF77;    16'd33187: out <= 16'h05AC;
    16'd33188: out <= 16'h034A;    16'd33189: out <= 16'h0421;    16'd33190: out <= 16'h00EC;    16'd33191: out <= 16'h0407;
    16'd33192: out <= 16'h0627;    16'd33193: out <= 16'h06A1;    16'd33194: out <= 16'hFEDB;    16'd33195: out <= 16'h0161;
    16'd33196: out <= 16'hFFE7;    16'd33197: out <= 16'hFE50;    16'd33198: out <= 16'h03DA;    16'd33199: out <= 16'h029D;
    16'd33200: out <= 16'h01D7;    16'd33201: out <= 16'h02E2;    16'd33202: out <= 16'h07DB;    16'd33203: out <= 16'h041E;
    16'd33204: out <= 16'h036C;    16'd33205: out <= 16'h0009;    16'd33206: out <= 16'h03CA;    16'd33207: out <= 16'h031D;
    16'd33208: out <= 16'h0375;    16'd33209: out <= 16'h0560;    16'd33210: out <= 16'h06CD;    16'd33211: out <= 16'hFEFB;
    16'd33212: out <= 16'h07C0;    16'd33213: out <= 16'h003E;    16'd33214: out <= 16'h0894;    16'd33215: out <= 16'h079B;
    16'd33216: out <= 16'hFE90;    16'd33217: out <= 16'h001B;    16'd33218: out <= 16'h018C;    16'd33219: out <= 16'h050A;
    16'd33220: out <= 16'h0520;    16'd33221: out <= 16'h02B5;    16'd33222: out <= 16'h019C;    16'd33223: out <= 16'h0BF6;
    16'd33224: out <= 16'h06DF;    16'd33225: out <= 16'h02C5;    16'd33226: out <= 16'h04F2;    16'd33227: out <= 16'h013C;
    16'd33228: out <= 16'h0544;    16'd33229: out <= 16'h0860;    16'd33230: out <= 16'h013F;    16'd33231: out <= 16'h0649;
    16'd33232: out <= 16'h04A7;    16'd33233: out <= 16'h0171;    16'd33234: out <= 16'hFE10;    16'd33235: out <= 16'h01D1;
    16'd33236: out <= 16'h08A9;    16'd33237: out <= 16'h0362;    16'd33238: out <= 16'h0829;    16'd33239: out <= 16'h0327;
    16'd33240: out <= 16'h077D;    16'd33241: out <= 16'h0247;    16'd33242: out <= 16'hFDE0;    16'd33243: out <= 16'h0111;
    16'd33244: out <= 16'h0111;    16'd33245: out <= 16'h0415;    16'd33246: out <= 16'h075B;    16'd33247: out <= 16'hFE08;
    16'd33248: out <= 16'h0320;    16'd33249: out <= 16'h09F9;    16'd33250: out <= 16'h056C;    16'd33251: out <= 16'h0699;
    16'd33252: out <= 16'h03C2;    16'd33253: out <= 16'hFD98;    16'd33254: out <= 16'h07A3;    16'd33255: out <= 16'hFC77;
    16'd33256: out <= 16'h00B3;    16'd33257: out <= 16'hFEB2;    16'd33258: out <= 16'h07B1;    16'd33259: out <= 16'h0038;
    16'd33260: out <= 16'h049C;    16'd33261: out <= 16'h032F;    16'd33262: out <= 16'hFF93;    16'd33263: out <= 16'hFF2B;
    16'd33264: out <= 16'h031D;    16'd33265: out <= 16'h000C;    16'd33266: out <= 16'h017D;    16'd33267: out <= 16'hFB80;
    16'd33268: out <= 16'hFADD;    16'd33269: out <= 16'hFC89;    16'd33270: out <= 16'hFBD9;    16'd33271: out <= 16'h0212;
    16'd33272: out <= 16'hFCD1;    16'd33273: out <= 16'h073E;    16'd33274: out <= 16'hFEFA;    16'd33275: out <= 16'h0503;
    16'd33276: out <= 16'h0484;    16'd33277: out <= 16'h00F2;    16'd33278: out <= 16'h0283;    16'd33279: out <= 16'h007E;
    16'd33280: out <= 16'h05D8;    16'd33281: out <= 16'hFE4D;    16'd33282: out <= 16'h0202;    16'd33283: out <= 16'h033D;
    16'd33284: out <= 16'h0084;    16'd33285: out <= 16'h0056;    16'd33286: out <= 16'hFAE7;    16'd33287: out <= 16'hFCCE;
    16'd33288: out <= 16'hFA46;    16'd33289: out <= 16'hFBBB;    16'd33290: out <= 16'h03F6;    16'd33291: out <= 16'h00B3;
    16'd33292: out <= 16'hFF24;    16'd33293: out <= 16'h0079;    16'd33294: out <= 16'hFF10;    16'd33295: out <= 16'h0186;
    16'd33296: out <= 16'hFE04;    16'd33297: out <= 16'h033C;    16'd33298: out <= 16'h03DA;    16'd33299: out <= 16'hFDBB;
    16'd33300: out <= 16'hFCFF;    16'd33301: out <= 16'h01C3;    16'd33302: out <= 16'h0512;    16'd33303: out <= 16'h0442;
    16'd33304: out <= 16'h05D0;    16'd33305: out <= 16'h06A6;    16'd33306: out <= 16'h002A;    16'd33307: out <= 16'h0332;
    16'd33308: out <= 16'hFFA7;    16'd33309: out <= 16'h00DB;    16'd33310: out <= 16'h0371;    16'd33311: out <= 16'hFE82;
    16'd33312: out <= 16'h0260;    16'd33313: out <= 16'h01BC;    16'd33314: out <= 16'h087C;    16'd33315: out <= 16'h07CC;
    16'd33316: out <= 16'h04C6;    16'd33317: out <= 16'h0042;    16'd33318: out <= 16'h03A5;    16'd33319: out <= 16'h03CB;
    16'd33320: out <= 16'hFFE5;    16'd33321: out <= 16'h078C;    16'd33322: out <= 16'h08DA;    16'd33323: out <= 16'h00A2;
    16'd33324: out <= 16'h07CA;    16'd33325: out <= 16'h04E1;    16'd33326: out <= 16'h04BA;    16'd33327: out <= 16'hFE3B;
    16'd33328: out <= 16'h0AA0;    16'd33329: out <= 16'h0460;    16'd33330: out <= 16'hFB95;    16'd33331: out <= 16'h06C3;
    16'd33332: out <= 16'hFED3;    16'd33333: out <= 16'h0691;    16'd33334: out <= 16'h0110;    16'd33335: out <= 16'h016F;
    16'd33336: out <= 16'h0717;    16'd33337: out <= 16'h0696;    16'd33338: out <= 16'hFC10;    16'd33339: out <= 16'hFF26;
    16'd33340: out <= 16'h0451;    16'd33341: out <= 16'h0551;    16'd33342: out <= 16'h095D;    16'd33343: out <= 16'h06AB;
    16'd33344: out <= 16'h01BF;    16'd33345: out <= 16'h04E5;    16'd33346: out <= 16'h022B;    16'd33347: out <= 16'h00A9;
    16'd33348: out <= 16'h04F9;    16'd33349: out <= 16'h07F1;    16'd33350: out <= 16'h093F;    16'd33351: out <= 16'h055B;
    16'd33352: out <= 16'h0E03;    16'd33353: out <= 16'h0B2E;    16'd33354: out <= 16'h05DE;    16'd33355: out <= 16'h0113;
    16'd33356: out <= 16'h05BE;    16'd33357: out <= 16'h04BD;    16'd33358: out <= 16'h05E3;    16'd33359: out <= 16'h0779;
    16'd33360: out <= 16'h0130;    16'd33361: out <= 16'h0253;    16'd33362: out <= 16'h0290;    16'd33363: out <= 16'h039D;
    16'd33364: out <= 16'h03C5;    16'd33365: out <= 16'h071E;    16'd33366: out <= 16'h0A00;    16'd33367: out <= 16'h0256;
    16'd33368: out <= 16'h0220;    16'd33369: out <= 16'h0891;    16'd33370: out <= 16'h025C;    16'd33371: out <= 16'hFFA1;
    16'd33372: out <= 16'h0205;    16'd33373: out <= 16'h076D;    16'd33374: out <= 16'h03D8;    16'd33375: out <= 16'h03B8;
    16'd33376: out <= 16'hFA0D;    16'd33377: out <= 16'h0275;    16'd33378: out <= 16'h07E2;    16'd33379: out <= 16'h055A;
    16'd33380: out <= 16'h0621;    16'd33381: out <= 16'h0623;    16'd33382: out <= 16'h0759;    16'd33383: out <= 16'h0757;
    16'd33384: out <= 16'h03F9;    16'd33385: out <= 16'h0B25;    16'd33386: out <= 16'h0A3D;    16'd33387: out <= 16'h03E2;
    16'd33388: out <= 16'hFFF9;    16'd33389: out <= 16'hFCCD;    16'd33390: out <= 16'h040C;    16'd33391: out <= 16'hFB5C;
    16'd33392: out <= 16'hFE6E;    16'd33393: out <= 16'h024E;    16'd33394: out <= 16'hFFBD;    16'd33395: out <= 16'h0593;
    16'd33396: out <= 16'h014F;    16'd33397: out <= 16'h0486;    16'd33398: out <= 16'hFFAA;    16'd33399: out <= 16'h0416;
    16'd33400: out <= 16'h06FB;    16'd33401: out <= 16'h042C;    16'd33402: out <= 16'h03BD;    16'd33403: out <= 16'h05AD;
    16'd33404: out <= 16'h047E;    16'd33405: out <= 16'h0A72;    16'd33406: out <= 16'h02B6;    16'd33407: out <= 16'hFF03;
    16'd33408: out <= 16'h051F;    16'd33409: out <= 16'h047A;    16'd33410: out <= 16'h0458;    16'd33411: out <= 16'h05ED;
    16'd33412: out <= 16'h00EF;    16'd33413: out <= 16'h02F1;    16'd33414: out <= 16'h065A;    16'd33415: out <= 16'h06B1;
    16'd33416: out <= 16'hFF2D;    16'd33417: out <= 16'h0460;    16'd33418: out <= 16'h05C6;    16'd33419: out <= 16'h04C9;
    16'd33420: out <= 16'h04CF;    16'd33421: out <= 16'hFF8B;    16'd33422: out <= 16'h04E4;    16'd33423: out <= 16'h0BF9;
    16'd33424: out <= 16'hFBC0;    16'd33425: out <= 16'h0097;    16'd33426: out <= 16'h0215;    16'd33427: out <= 16'h0488;
    16'd33428: out <= 16'h0452;    16'd33429: out <= 16'h01CB;    16'd33430: out <= 16'h032B;    16'd33431: out <= 16'h0141;
    16'd33432: out <= 16'h0FCC;    16'd33433: out <= 16'h03CB;    16'd33434: out <= 16'h0462;    16'd33435: out <= 16'h0003;
    16'd33436: out <= 16'h0836;    16'd33437: out <= 16'h0783;    16'd33438: out <= 16'h006C;    16'd33439: out <= 16'h0198;
    16'd33440: out <= 16'h03DE;    16'd33441: out <= 16'h04DE;    16'd33442: out <= 16'h02FD;    16'd33443: out <= 16'hFF6F;
    16'd33444: out <= 16'h0708;    16'd33445: out <= 16'hFF4C;    16'd33446: out <= 16'h0432;    16'd33447: out <= 16'h062B;
    16'd33448: out <= 16'hFFB3;    16'd33449: out <= 16'h0A58;    16'd33450: out <= 16'h07D1;    16'd33451: out <= 16'h0A4F;
    16'd33452: out <= 16'h05CA;    16'd33453: out <= 16'hFC90;    16'd33454: out <= 16'h05C8;    16'd33455: out <= 16'h0728;
    16'd33456: out <= 16'h076B;    16'd33457: out <= 16'h09E1;    16'd33458: out <= 16'h093F;    16'd33459: out <= 16'h00CD;
    16'd33460: out <= 16'h020D;    16'd33461: out <= 16'h0CC4;    16'd33462: out <= 16'h024F;    16'd33463: out <= 16'h020C;
    16'd33464: out <= 16'h08B8;    16'd33465: out <= 16'h0072;    16'd33466: out <= 16'hFEC4;    16'd33467: out <= 16'h0575;
    16'd33468: out <= 16'h04FD;    16'd33469: out <= 16'h0198;    16'd33470: out <= 16'h077A;    16'd33471: out <= 16'h0853;
    16'd33472: out <= 16'h0725;    16'd33473: out <= 16'h0B9D;    16'd33474: out <= 16'hFD92;    16'd33475: out <= 16'h0493;
    16'd33476: out <= 16'hFEAA;    16'd33477: out <= 16'hFB6D;    16'd33478: out <= 16'h05D6;    16'd33479: out <= 16'h070B;
    16'd33480: out <= 16'hFF86;    16'd33481: out <= 16'h067A;    16'd33482: out <= 16'h00A7;    16'd33483: out <= 16'h05AA;
    16'd33484: out <= 16'h047B;    16'd33485: out <= 16'h0084;    16'd33486: out <= 16'hFCD4;    16'd33487: out <= 16'h0491;
    16'd33488: out <= 16'h0125;    16'd33489: out <= 16'h0103;    16'd33490: out <= 16'h08CC;    16'd33491: out <= 16'h038F;
    16'd33492: out <= 16'h00B4;    16'd33493: out <= 16'h0882;    16'd33494: out <= 16'h004D;    16'd33495: out <= 16'h04CB;
    16'd33496: out <= 16'h03D9;    16'd33497: out <= 16'h030A;    16'd33498: out <= 16'h0266;    16'd33499: out <= 16'h0609;
    16'd33500: out <= 16'h01E3;    16'd33501: out <= 16'h0841;    16'd33502: out <= 16'h00DE;    16'd33503: out <= 16'h0299;
    16'd33504: out <= 16'h03A1;    16'd33505: out <= 16'h038E;    16'd33506: out <= 16'h058B;    16'd33507: out <= 16'h0026;
    16'd33508: out <= 16'h0207;    16'd33509: out <= 16'h058D;    16'd33510: out <= 16'h0311;    16'd33511: out <= 16'hFE68;
    16'd33512: out <= 16'hFEF7;    16'd33513: out <= 16'hF9BE;    16'd33514: out <= 16'hF6EC;    16'd33515: out <= 16'hFDF9;
    16'd33516: out <= 16'hFF4B;    16'd33517: out <= 16'h0141;    16'd33518: out <= 16'h0189;    16'd33519: out <= 16'hFE66;
    16'd33520: out <= 16'hFFE9;    16'd33521: out <= 16'hFBC4;    16'd33522: out <= 16'h020D;    16'd33523: out <= 16'h00A2;
    16'd33524: out <= 16'h0077;    16'd33525: out <= 16'hFCFB;    16'd33526: out <= 16'hFD87;    16'd33527: out <= 16'hFF0A;
    16'd33528: out <= 16'h048F;    16'd33529: out <= 16'hFE0B;    16'd33530: out <= 16'h00D3;    16'd33531: out <= 16'hFBD1;
    16'd33532: out <= 16'h0459;    16'd33533: out <= 16'h058D;    16'd33534: out <= 16'hFDA4;    16'd33535: out <= 16'h040E;
    16'd33536: out <= 16'h0357;    16'd33537: out <= 16'hFB32;    16'd33538: out <= 16'h0133;    16'd33539: out <= 16'hFFEC;
    16'd33540: out <= 16'h00A2;    16'd33541: out <= 16'h00F8;    16'd33542: out <= 16'hFE7C;    16'd33543: out <= 16'hF899;
    16'd33544: out <= 16'h0B8F;    16'd33545: out <= 16'h00A1;    16'd33546: out <= 16'h066D;    16'd33547: out <= 16'h0576;
    16'd33548: out <= 16'hF93C;    16'd33549: out <= 16'hF94A;    16'd33550: out <= 16'h0691;    16'd33551: out <= 16'hFE46;
    16'd33552: out <= 16'h0357;    16'd33553: out <= 16'h0117;    16'd33554: out <= 16'hFFD6;    16'd33555: out <= 16'hFDA8;
    16'd33556: out <= 16'h011E;    16'd33557: out <= 16'hFCA3;    16'd33558: out <= 16'h0021;    16'd33559: out <= 16'h0112;
    16'd33560: out <= 16'h04FC;    16'd33561: out <= 16'h0564;    16'd33562: out <= 16'h0277;    16'd33563: out <= 16'h0735;
    16'd33564: out <= 16'hFD34;    16'd33565: out <= 16'h04BC;    16'd33566: out <= 16'h070F;    16'd33567: out <= 16'h0875;
    16'd33568: out <= 16'h0888;    16'd33569: out <= 16'h0AEF;    16'd33570: out <= 16'hFE86;    16'd33571: out <= 16'hFBFA;
    16'd33572: out <= 16'h0398;    16'd33573: out <= 16'h020D;    16'd33574: out <= 16'h04F8;    16'd33575: out <= 16'h02B7;
    16'd33576: out <= 16'h07AD;    16'd33577: out <= 16'h028A;    16'd33578: out <= 16'h0415;    16'd33579: out <= 16'h0AA8;
    16'd33580: out <= 16'hFF7D;    16'd33581: out <= 16'h058C;    16'd33582: out <= 16'h05F0;    16'd33583: out <= 16'hFE6B;
    16'd33584: out <= 16'h060C;    16'd33585: out <= 16'h04E6;    16'd33586: out <= 16'h0687;    16'd33587: out <= 16'h02A0;
    16'd33588: out <= 16'h01FC;    16'd33589: out <= 16'h03DA;    16'd33590: out <= 16'h0215;    16'd33591: out <= 16'h048B;
    16'd33592: out <= 16'hFEC0;    16'd33593: out <= 16'h02A0;    16'd33594: out <= 16'h065F;    16'd33595: out <= 16'h057E;
    16'd33596: out <= 16'h0A75;    16'd33597: out <= 16'h05C8;    16'd33598: out <= 16'h0236;    16'd33599: out <= 16'h0444;
    16'd33600: out <= 16'hFDB2;    16'd33601: out <= 16'hFF87;    16'd33602: out <= 16'h0945;    16'd33603: out <= 16'h04A8;
    16'd33604: out <= 16'h02E3;    16'd33605: out <= 16'h06EE;    16'd33606: out <= 16'h01F0;    16'd33607: out <= 16'h02E8;
    16'd33608: out <= 16'h004E;    16'd33609: out <= 16'h0D52;    16'd33610: out <= 16'hFCE2;    16'd33611: out <= 16'h055C;
    16'd33612: out <= 16'h08EE;    16'd33613: out <= 16'h07A6;    16'd33614: out <= 16'h0487;    16'd33615: out <= 16'h0B57;
    16'd33616: out <= 16'h02A8;    16'd33617: out <= 16'h0750;    16'd33618: out <= 16'h0538;    16'd33619: out <= 16'h095D;
    16'd33620: out <= 16'h0784;    16'd33621: out <= 16'h04A9;    16'd33622: out <= 16'h0708;    16'd33623: out <= 16'h023D;
    16'd33624: out <= 16'hFBED;    16'd33625: out <= 16'h0AA3;    16'd33626: out <= 16'hFF49;    16'd33627: out <= 16'h0020;
    16'd33628: out <= 16'hFEC0;    16'd33629: out <= 16'h067A;    16'd33630: out <= 16'h00B2;    16'd33631: out <= 16'h08A9;
    16'd33632: out <= 16'h0417;    16'd33633: out <= 16'h016C;    16'd33634: out <= 16'hFDEF;    16'd33635: out <= 16'h08CE;
    16'd33636: out <= 16'h039F;    16'd33637: out <= 16'h056D;    16'd33638: out <= 16'h04CB;    16'd33639: out <= 16'h0276;
    16'd33640: out <= 16'h09A9;    16'd33641: out <= 16'hFE78;    16'd33642: out <= 16'h0303;    16'd33643: out <= 16'h0CB6;
    16'd33644: out <= 16'hFE70;    16'd33645: out <= 16'h03E6;    16'd33646: out <= 16'h07E8;    16'd33647: out <= 16'h04FB;
    16'd33648: out <= 16'h00D0;    16'd33649: out <= 16'h071E;    16'd33650: out <= 16'h08B8;    16'd33651: out <= 16'hFFD5;
    16'd33652: out <= 16'h0415;    16'd33653: out <= 16'h05B3;    16'd33654: out <= 16'h0578;    16'd33655: out <= 16'h0061;
    16'd33656: out <= 16'h04E0;    16'd33657: out <= 16'h0452;    16'd33658: out <= 16'h06EA;    16'd33659: out <= 16'h0569;
    16'd33660: out <= 16'h0E4D;    16'd33661: out <= 16'h05F5;    16'd33662: out <= 16'h04B1;    16'd33663: out <= 16'h062A;
    16'd33664: out <= 16'h03D6;    16'd33665: out <= 16'h0B0D;    16'd33666: out <= 16'h0531;    16'd33667: out <= 16'h0B40;
    16'd33668: out <= 16'h04A3;    16'd33669: out <= 16'h035F;    16'd33670: out <= 16'h0386;    16'd33671: out <= 16'h0348;
    16'd33672: out <= 16'h0A0B;    16'd33673: out <= 16'h01D6;    16'd33674: out <= 16'h04F4;    16'd33675: out <= 16'h03B4;
    16'd33676: out <= 16'h04BB;    16'd33677: out <= 16'h04A4;    16'd33678: out <= 16'hFF3E;    16'd33679: out <= 16'h0312;
    16'd33680: out <= 16'h06A8;    16'd33681: out <= 16'h014E;    16'd33682: out <= 16'h0650;    16'd33683: out <= 16'hFD3F;
    16'd33684: out <= 16'h04DB;    16'd33685: out <= 16'h0386;    16'd33686: out <= 16'h04F0;    16'd33687: out <= 16'h02FC;
    16'd33688: out <= 16'h0234;    16'd33689: out <= 16'h079A;    16'd33690: out <= 16'h03DA;    16'd33691: out <= 16'h054F;
    16'd33692: out <= 16'h097F;    16'd33693: out <= 16'h0913;    16'd33694: out <= 16'h060C;    16'd33695: out <= 16'h03BC;
    16'd33696: out <= 16'h01E9;    16'd33697: out <= 16'h0074;    16'd33698: out <= 16'h053C;    16'd33699: out <= 16'h04AD;
    16'd33700: out <= 16'hFFA6;    16'd33701: out <= 16'hFC35;    16'd33702: out <= 16'h0724;    16'd33703: out <= 16'h09A4;
    16'd33704: out <= 16'h078C;    16'd33705: out <= 16'h01AF;    16'd33706: out <= 16'hF7C9;    16'd33707: out <= 16'h05D3;
    16'd33708: out <= 16'hFF90;    16'd33709: out <= 16'h0694;    16'd33710: out <= 16'h0573;    16'd33711: out <= 16'h0239;
    16'd33712: out <= 16'h0854;    16'd33713: out <= 16'h078F;    16'd33714: out <= 16'h02B7;    16'd33715: out <= 16'h0A5F;
    16'd33716: out <= 16'h011F;    16'd33717: out <= 16'h0161;    16'd33718: out <= 16'h0696;    16'd33719: out <= 16'h036B;
    16'd33720: out <= 16'hFE06;    16'd33721: out <= 16'h0606;    16'd33722: out <= 16'h06F7;    16'd33723: out <= 16'hFC57;
    16'd33724: out <= 16'h03ED;    16'd33725: out <= 16'h0446;    16'd33726: out <= 16'hFEC3;    16'd33727: out <= 16'h0C48;
    16'd33728: out <= 16'hFF9F;    16'd33729: out <= 16'h0217;    16'd33730: out <= 16'h04B4;    16'd33731: out <= 16'h027F;
    16'd33732: out <= 16'h0769;    16'd33733: out <= 16'h0692;    16'd33734: out <= 16'h0241;    16'd33735: out <= 16'h053F;
    16'd33736: out <= 16'hFFCE;    16'd33737: out <= 16'hFED7;    16'd33738: out <= 16'h006D;    16'd33739: out <= 16'hFF0D;
    16'd33740: out <= 16'h0034;    16'd33741: out <= 16'h0289;    16'd33742: out <= 16'h07D2;    16'd33743: out <= 16'h0978;
    16'd33744: out <= 16'h0675;    16'd33745: out <= 16'h05C5;    16'd33746: out <= 16'h0154;    16'd33747: out <= 16'h06E3;
    16'd33748: out <= 16'h00C8;    16'd33749: out <= 16'h0928;    16'd33750: out <= 16'h0974;    16'd33751: out <= 16'h077F;
    16'd33752: out <= 16'h06AE;    16'd33753: out <= 16'hFFD0;    16'd33754: out <= 16'h01BB;    16'd33755: out <= 16'h049E;
    16'd33756: out <= 16'hFEB4;    16'd33757: out <= 16'h0860;    16'd33758: out <= 16'h05BC;    16'd33759: out <= 16'h0560;
    16'd33760: out <= 16'h03A6;    16'd33761: out <= 16'h05F5;    16'd33762: out <= 16'h06E9;    16'd33763: out <= 16'h023B;
    16'd33764: out <= 16'h0995;    16'd33765: out <= 16'hFAD7;    16'd33766: out <= 16'h046A;    16'd33767: out <= 16'h025A;
    16'd33768: out <= 16'h04E3;    16'd33769: out <= 16'h0264;    16'd33770: out <= 16'h00B2;    16'd33771: out <= 16'h002D;
    16'd33772: out <= 16'h01C2;    16'd33773: out <= 16'h005B;    16'd33774: out <= 16'h0026;    16'd33775: out <= 16'h05F2;
    16'd33776: out <= 16'hFA61;    16'd33777: out <= 16'hFED9;    16'd33778: out <= 16'h02EA;    16'd33779: out <= 16'h03E3;
    16'd33780: out <= 16'h0201;    16'd33781: out <= 16'h07A8;    16'd33782: out <= 16'hFF5F;    16'd33783: out <= 16'hFBF3;
    16'd33784: out <= 16'hFFF5;    16'd33785: out <= 16'h03BA;    16'd33786: out <= 16'h0085;    16'd33787: out <= 16'hFFA6;
    16'd33788: out <= 16'hFDD2;    16'd33789: out <= 16'h0000;    16'd33790: out <= 16'hFBB4;    16'd33791: out <= 16'h037D;
    16'd33792: out <= 16'hFB98;    16'd33793: out <= 16'hFF41;    16'd33794: out <= 16'hFDF1;    16'd33795: out <= 16'hFE75;
    16'd33796: out <= 16'hFB75;    16'd33797: out <= 16'h03B5;    16'd33798: out <= 16'hF811;    16'd33799: out <= 16'hFD87;
    16'd33800: out <= 16'hFE6D;    16'd33801: out <= 16'hFB64;    16'd33802: out <= 16'hFE58;    16'd33803: out <= 16'hF8D7;
    16'd33804: out <= 16'hFE0A;    16'd33805: out <= 16'hFE4A;    16'd33806: out <= 16'hFD37;    16'd33807: out <= 16'h0452;
    16'd33808: out <= 16'h029A;    16'd33809: out <= 16'h0460;    16'd33810: out <= 16'h072A;    16'd33811: out <= 16'h0381;
    16'd33812: out <= 16'h0096;    16'd33813: out <= 16'hFA63;    16'd33814: out <= 16'hF8DC;    16'd33815: out <= 16'h058B;
    16'd33816: out <= 16'h0135;    16'd33817: out <= 16'h034E;    16'd33818: out <= 16'h0138;    16'd33819: out <= 16'h01DB;
    16'd33820: out <= 16'h027C;    16'd33821: out <= 16'h0454;    16'd33822: out <= 16'h03EB;    16'd33823: out <= 16'h0453;
    16'd33824: out <= 16'h027B;    16'd33825: out <= 16'h059E;    16'd33826: out <= 16'h0359;    16'd33827: out <= 16'h06D2;
    16'd33828: out <= 16'h07EC;    16'd33829: out <= 16'h09EB;    16'd33830: out <= 16'h00A2;    16'd33831: out <= 16'h0055;
    16'd33832: out <= 16'h083C;    16'd33833: out <= 16'h0198;    16'd33834: out <= 16'hFF07;    16'd33835: out <= 16'h031E;
    16'd33836: out <= 16'h0598;    16'd33837: out <= 16'h0314;    16'd33838: out <= 16'h0496;    16'd33839: out <= 16'h0934;
    16'd33840: out <= 16'h0727;    16'd33841: out <= 16'h02B4;    16'd33842: out <= 16'hFD21;    16'd33843: out <= 16'h0372;
    16'd33844: out <= 16'h05B1;    16'd33845: out <= 16'h06FF;    16'd33846: out <= 16'hFB1D;    16'd33847: out <= 16'h03FB;
    16'd33848: out <= 16'h040D;    16'd33849: out <= 16'h059F;    16'd33850: out <= 16'h0000;    16'd33851: out <= 16'h04C4;
    16'd33852: out <= 16'h0893;    16'd33853: out <= 16'hFDE2;    16'd33854: out <= 16'h0194;    16'd33855: out <= 16'h09E0;
    16'd33856: out <= 16'h0258;    16'd33857: out <= 16'h05BB;    16'd33858: out <= 16'h06E0;    16'd33859: out <= 16'h0319;
    16'd33860: out <= 16'h0047;    16'd33861: out <= 16'h0670;    16'd33862: out <= 16'h0654;    16'd33863: out <= 16'hFEA1;
    16'd33864: out <= 16'h0784;    16'd33865: out <= 16'h0462;    16'd33866: out <= 16'hFFE0;    16'd33867: out <= 16'h0706;
    16'd33868: out <= 16'h055C;    16'd33869: out <= 16'h019E;    16'd33870: out <= 16'h0277;    16'd33871: out <= 16'h02F1;
    16'd33872: out <= 16'h03D5;    16'd33873: out <= 16'h02FA;    16'd33874: out <= 16'hFE08;    16'd33875: out <= 16'h00AE;
    16'd33876: out <= 16'h0C33;    16'd33877: out <= 16'h075B;    16'd33878: out <= 16'hFBC0;    16'd33879: out <= 16'h0C0B;
    16'd33880: out <= 16'h02B3;    16'd33881: out <= 16'h05E0;    16'd33882: out <= 16'h050A;    16'd33883: out <= 16'h0566;
    16'd33884: out <= 16'h0147;    16'd33885: out <= 16'hFF36;    16'd33886: out <= 16'h02B1;    16'd33887: out <= 16'h05BE;
    16'd33888: out <= 16'h049B;    16'd33889: out <= 16'h0349;    16'd33890: out <= 16'h02E7;    16'd33891: out <= 16'h0496;
    16'd33892: out <= 16'h05B8;    16'd33893: out <= 16'hFF4D;    16'd33894: out <= 16'h00A9;    16'd33895: out <= 16'hFFCC;
    16'd33896: out <= 16'h062F;    16'd33897: out <= 16'hFBF5;    16'd33898: out <= 16'h0004;    16'd33899: out <= 16'h0286;
    16'd33900: out <= 16'h01DE;    16'd33901: out <= 16'h029F;    16'd33902: out <= 16'hFFD0;    16'd33903: out <= 16'h091D;
    16'd33904: out <= 16'h0ADD;    16'd33905: out <= 16'h06CA;    16'd33906: out <= 16'h04A1;    16'd33907: out <= 16'h06F0;
    16'd33908: out <= 16'h045B;    16'd33909: out <= 16'h05D0;    16'd33910: out <= 16'h044E;    16'd33911: out <= 16'h0930;
    16'd33912: out <= 16'h0530;    16'd33913: out <= 16'h0C85;    16'd33914: out <= 16'h0122;    16'd33915: out <= 16'h057C;
    16'd33916: out <= 16'h0E46;    16'd33917: out <= 16'hFF83;    16'd33918: out <= 16'h0EA1;    16'd33919: out <= 16'h0337;
    16'd33920: out <= 16'hF94B;    16'd33921: out <= 16'h08E5;    16'd33922: out <= 16'hFDC6;    16'd33923: out <= 16'h01E9;
    16'd33924: out <= 16'h0457;    16'd33925: out <= 16'h01CE;    16'd33926: out <= 16'h00D4;    16'd33927: out <= 16'h095A;
    16'd33928: out <= 16'hFBEA;    16'd33929: out <= 16'h06F3;    16'd33930: out <= 16'hFBB7;    16'd33931: out <= 16'h0079;
    16'd33932: out <= 16'h089A;    16'd33933: out <= 16'h026F;    16'd33934: out <= 16'h016C;    16'd33935: out <= 16'h02E0;
    16'd33936: out <= 16'hFFEF;    16'd33937: out <= 16'h0505;    16'd33938: out <= 16'h012E;    16'd33939: out <= 16'hFED9;
    16'd33940: out <= 16'h083B;    16'd33941: out <= 16'hFB33;    16'd33942: out <= 16'h041E;    16'd33943: out <= 16'h01B2;
    16'd33944: out <= 16'h098C;    16'd33945: out <= 16'h0528;    16'd33946: out <= 16'h0346;    16'd33947: out <= 16'hFF94;
    16'd33948: out <= 16'h0C48;    16'd33949: out <= 16'hFEB6;    16'd33950: out <= 16'hFF5D;    16'd33951: out <= 16'h00EF;
    16'd33952: out <= 16'h060B;    16'd33953: out <= 16'h0574;    16'd33954: out <= 16'hFB88;    16'd33955: out <= 16'h01E7;
    16'd33956: out <= 16'h033D;    16'd33957: out <= 16'hFF95;    16'd33958: out <= 16'h0658;    16'd33959: out <= 16'h08B0;
    16'd33960: out <= 16'h0023;    16'd33961: out <= 16'h066E;    16'd33962: out <= 16'h065F;    16'd33963: out <= 16'h069A;
    16'd33964: out <= 16'h010E;    16'd33965: out <= 16'h0ACA;    16'd33966: out <= 16'h02F4;    16'd33967: out <= 16'h0A83;
    16'd33968: out <= 16'h090D;    16'd33969: out <= 16'h0027;    16'd33970: out <= 16'h000C;    16'd33971: out <= 16'hFF9D;
    16'd33972: out <= 16'h04ED;    16'd33973: out <= 16'hFBEA;    16'd33974: out <= 16'h06AA;    16'd33975: out <= 16'h0A38;
    16'd33976: out <= 16'h04F3;    16'd33977: out <= 16'h0737;    16'd33978: out <= 16'h04FF;    16'd33979: out <= 16'h064E;
    16'd33980: out <= 16'h0345;    16'd33981: out <= 16'hFE9A;    16'd33982: out <= 16'h07A1;    16'd33983: out <= 16'h068B;
    16'd33984: out <= 16'h06AA;    16'd33985: out <= 16'h01B3;    16'd33986: out <= 16'h009B;    16'd33987: out <= 16'hFE7F;
    16'd33988: out <= 16'h037D;    16'd33989: out <= 16'h0999;    16'd33990: out <= 16'hFEA5;    16'd33991: out <= 16'h02CC;
    16'd33992: out <= 16'h000D;    16'd33993: out <= 16'h0518;    16'd33994: out <= 16'h07AB;    16'd33995: out <= 16'h063B;
    16'd33996: out <= 16'hFEDB;    16'd33997: out <= 16'h01D0;    16'd33998: out <= 16'h08D5;    16'd33999: out <= 16'h0741;
    16'd34000: out <= 16'h046E;    16'd34001: out <= 16'h00B3;    16'd34002: out <= 16'h094C;    16'd34003: out <= 16'h005E;
    16'd34004: out <= 16'h077D;    16'd34005: out <= 16'h0484;    16'd34006: out <= 16'h0642;    16'd34007: out <= 16'h0AA1;
    16'd34008: out <= 16'h022F;    16'd34009: out <= 16'hFF9D;    16'd34010: out <= 16'h0740;    16'd34011: out <= 16'hFF4D;
    16'd34012: out <= 16'h01E3;    16'd34013: out <= 16'h0638;    16'd34014: out <= 16'h0519;    16'd34015: out <= 16'h05C9;
    16'd34016: out <= 16'h0278;    16'd34017: out <= 16'h06BE;    16'd34018: out <= 16'h01FF;    16'd34019: out <= 16'h03F1;
    16'd34020: out <= 16'h02AA;    16'd34021: out <= 16'h095B;    16'd34022: out <= 16'h024D;    16'd34023: out <= 16'hFF34;
    16'd34024: out <= 16'h0234;    16'd34025: out <= 16'h06B1;    16'd34026: out <= 16'h0572;    16'd34027: out <= 16'h04FA;
    16'd34028: out <= 16'h02ED;    16'd34029: out <= 16'hF7F4;    16'd34030: out <= 16'hFF83;    16'd34031: out <= 16'h0045;
    16'd34032: out <= 16'h00A0;    16'd34033: out <= 16'h081B;    16'd34034: out <= 16'h0525;    16'd34035: out <= 16'hFEAB;
    16'd34036: out <= 16'h0282;    16'd34037: out <= 16'hFC21;    16'd34038: out <= 16'hFBD7;    16'd34039: out <= 16'hFF2B;
    16'd34040: out <= 16'h00B5;    16'd34041: out <= 16'hFFA8;    16'd34042: out <= 16'hFFDC;    16'd34043: out <= 16'hFF66;
    16'd34044: out <= 16'h02B8;    16'd34045: out <= 16'hFFEF;    16'd34046: out <= 16'hFC94;    16'd34047: out <= 16'hFBE3;
    16'd34048: out <= 16'h0002;    16'd34049: out <= 16'hFCF1;    16'd34050: out <= 16'h01D8;    16'd34051: out <= 16'hFFAC;
    16'd34052: out <= 16'h04D3;    16'd34053: out <= 16'hFBC2;    16'd34054: out <= 16'hFB53;    16'd34055: out <= 16'hFE4C;
    16'd34056: out <= 16'h030B;    16'd34057: out <= 16'h01B8;    16'd34058: out <= 16'hFCA7;    16'd34059: out <= 16'h01CF;
    16'd34060: out <= 16'h01CB;    16'd34061: out <= 16'hFB14;    16'd34062: out <= 16'hFC98;    16'd34063: out <= 16'hFA1B;
    16'd34064: out <= 16'hFEB6;    16'd34065: out <= 16'hFAAD;    16'd34066: out <= 16'hFE0F;    16'd34067: out <= 16'h0416;
    16'd34068: out <= 16'h0019;    16'd34069: out <= 16'h056B;    16'd34070: out <= 16'h057E;    16'd34071: out <= 16'h076E;
    16'd34072: out <= 16'hFD7A;    16'd34073: out <= 16'h0117;    16'd34074: out <= 16'hFED7;    16'd34075: out <= 16'h0859;
    16'd34076: out <= 16'hF8B3;    16'd34077: out <= 16'h0169;    16'd34078: out <= 16'h0156;    16'd34079: out <= 16'h0020;
    16'd34080: out <= 16'h0660;    16'd34081: out <= 16'h0967;    16'd34082: out <= 16'h0193;    16'd34083: out <= 16'h030A;
    16'd34084: out <= 16'h098D;    16'd34085: out <= 16'h079C;    16'd34086: out <= 16'h075F;    16'd34087: out <= 16'h03F5;
    16'd34088: out <= 16'h01B4;    16'd34089: out <= 16'h05D1;    16'd34090: out <= 16'h059F;    16'd34091: out <= 16'hFE7B;
    16'd34092: out <= 16'h0A27;    16'd34093: out <= 16'h0387;    16'd34094: out <= 16'h035E;    16'd34095: out <= 16'hFF74;
    16'd34096: out <= 16'h0762;    16'd34097: out <= 16'h0B01;    16'd34098: out <= 16'h0127;    16'd34099: out <= 16'h030E;
    16'd34100: out <= 16'h04B5;    16'd34101: out <= 16'h08DC;    16'd34102: out <= 16'h0514;    16'd34103: out <= 16'h0DCA;
    16'd34104: out <= 16'h0576;    16'd34105: out <= 16'h057C;    16'd34106: out <= 16'h019F;    16'd34107: out <= 16'hFEEE;
    16'd34108: out <= 16'h043D;    16'd34109: out <= 16'h0936;    16'd34110: out <= 16'h052A;    16'd34111: out <= 16'h053D;
    16'd34112: out <= 16'h0224;    16'd34113: out <= 16'h04B4;    16'd34114: out <= 16'h01C0;    16'd34115: out <= 16'h085B;
    16'd34116: out <= 16'h04DA;    16'd34117: out <= 16'h0E0D;    16'd34118: out <= 16'h09C5;    16'd34119: out <= 16'h0ECF;
    16'd34120: out <= 16'h0192;    16'd34121: out <= 16'hFEE2;    16'd34122: out <= 16'h09C8;    16'd34123: out <= 16'h0378;
    16'd34124: out <= 16'h0A55;    16'd34125: out <= 16'hFFB7;    16'd34126: out <= 16'h0AAE;    16'd34127: out <= 16'h094F;
    16'd34128: out <= 16'hFE1C;    16'd34129: out <= 16'h08C9;    16'd34130: out <= 16'h026F;    16'd34131: out <= 16'h0580;
    16'd34132: out <= 16'h00E7;    16'd34133: out <= 16'hFFEE;    16'd34134: out <= 16'h06C7;    16'd34135: out <= 16'h0561;
    16'd34136: out <= 16'h0566;    16'd34137: out <= 16'hFED4;    16'd34138: out <= 16'h0192;    16'd34139: out <= 16'hFF0B;
    16'd34140: out <= 16'h02ED;    16'd34141: out <= 16'h074E;    16'd34142: out <= 16'h033C;    16'd34143: out <= 16'h057B;
    16'd34144: out <= 16'h0613;    16'd34145: out <= 16'h0E13;    16'd34146: out <= 16'hFF0A;    16'd34147: out <= 16'hFA75;
    16'd34148: out <= 16'h033A;    16'd34149: out <= 16'h053B;    16'd34150: out <= 16'h07E4;    16'd34151: out <= 16'h044E;
    16'd34152: out <= 16'h0A56;    16'd34153: out <= 16'h075A;    16'd34154: out <= 16'h08F2;    16'd34155: out <= 16'h0681;
    16'd34156: out <= 16'h085C;    16'd34157: out <= 16'h0158;    16'd34158: out <= 16'hF9DD;    16'd34159: out <= 16'h05EC;
    16'd34160: out <= 16'h01C7;    16'd34161: out <= 16'h0734;    16'd34162: out <= 16'hFE92;    16'd34163: out <= 16'h06AD;
    16'd34164: out <= 16'h055B;    16'd34165: out <= 16'h078F;    16'd34166: out <= 16'h067A;    16'd34167: out <= 16'hFFF8;
    16'd34168: out <= 16'hFA37;    16'd34169: out <= 16'h0763;    16'd34170: out <= 16'h0BCA;    16'd34171: out <= 16'h0284;
    16'd34172: out <= 16'h0187;    16'd34173: out <= 16'h0861;    16'd34174: out <= 16'h01B2;    16'd34175: out <= 16'h05E7;
    16'd34176: out <= 16'h075D;    16'd34177: out <= 16'h07F0;    16'd34178: out <= 16'h0736;    16'd34179: out <= 16'h086E;
    16'd34180: out <= 16'h0473;    16'd34181: out <= 16'h003E;    16'd34182: out <= 16'h02DD;    16'd34183: out <= 16'h0590;
    16'd34184: out <= 16'h01BE;    16'd34185: out <= 16'h09E6;    16'd34186: out <= 16'h02D7;    16'd34187: out <= 16'h061B;
    16'd34188: out <= 16'hFF9D;    16'd34189: out <= 16'h092E;    16'd34190: out <= 16'h01A3;    16'd34191: out <= 16'h00FA;
    16'd34192: out <= 16'h0561;    16'd34193: out <= 16'h0753;    16'd34194: out <= 16'h0513;    16'd34195: out <= 16'h02DC;
    16'd34196: out <= 16'h00A7;    16'd34197: out <= 16'hFACE;    16'd34198: out <= 16'h0357;    16'd34199: out <= 16'hFEE6;
    16'd34200: out <= 16'h0604;    16'd34201: out <= 16'h0484;    16'd34202: out <= 16'h062F;    16'd34203: out <= 16'h054B;
    16'd34204: out <= 16'h03FC;    16'd34205: out <= 16'h046D;    16'd34206: out <= 16'h0768;    16'd34207: out <= 16'h0339;
    16'd34208: out <= 16'h04D6;    16'd34209: out <= 16'h0B19;    16'd34210: out <= 16'hFF4D;    16'd34211: out <= 16'h0127;
    16'd34212: out <= 16'h013E;    16'd34213: out <= 16'h09B0;    16'd34214: out <= 16'h064E;    16'd34215: out <= 16'hFD56;
    16'd34216: out <= 16'h019A;    16'd34217: out <= 16'h025F;    16'd34218: out <= 16'h0CD6;    16'd34219: out <= 16'h0BB6;
    16'd34220: out <= 16'h025E;    16'd34221: out <= 16'h0186;    16'd34222: out <= 16'h0263;    16'd34223: out <= 16'h056E;
    16'd34224: out <= 16'h0389;    16'd34225: out <= 16'h014F;    16'd34226: out <= 16'h088C;    16'd34227: out <= 16'hFDB6;
    16'd34228: out <= 16'h0251;    16'd34229: out <= 16'h025B;    16'd34230: out <= 16'h03AA;    16'd34231: out <= 16'h0238;
    16'd34232: out <= 16'h0973;    16'd34233: out <= 16'h0506;    16'd34234: out <= 16'h039A;    16'd34235: out <= 16'h05BC;
    16'd34236: out <= 16'h0198;    16'd34237: out <= 16'h069B;    16'd34238: out <= 16'h0D7E;    16'd34239: out <= 16'h061B;
    16'd34240: out <= 16'hFEA5;    16'd34241: out <= 16'h00D9;    16'd34242: out <= 16'h0532;    16'd34243: out <= 16'hFF2C;
    16'd34244: out <= 16'hFFA1;    16'd34245: out <= 16'h05EF;    16'd34246: out <= 16'h086C;    16'd34247: out <= 16'h00F7;
    16'd34248: out <= 16'h0834;    16'd34249: out <= 16'hF935;    16'd34250: out <= 16'h05DB;    16'd34251: out <= 16'h03DB;
    16'd34252: out <= 16'h017C;    16'd34253: out <= 16'hFF64;    16'd34254: out <= 16'h05D4;    16'd34255: out <= 16'hFBB4;
    16'd34256: out <= 16'h00A3;    16'd34257: out <= 16'h0607;    16'd34258: out <= 16'h0BEB;    16'd34259: out <= 16'hFEC9;
    16'd34260: out <= 16'h02E4;    16'd34261: out <= 16'h092B;    16'd34262: out <= 16'h0590;    16'd34263: out <= 16'hFE47;
    16'd34264: out <= 16'h06A1;    16'd34265: out <= 16'h04E0;    16'd34266: out <= 16'hFF2B;    16'd34267: out <= 16'hFDDD;
    16'd34268: out <= 16'h06D5;    16'd34269: out <= 16'h03CF;    16'd34270: out <= 16'h0403;    16'd34271: out <= 16'hFDD8;
    16'd34272: out <= 16'h05E2;    16'd34273: out <= 16'h046A;    16'd34274: out <= 16'h0468;    16'd34275: out <= 16'h05CE;
    16'd34276: out <= 16'hFCA9;    16'd34277: out <= 16'h030F;    16'd34278: out <= 16'h03A9;    16'd34279: out <= 16'h01C3;
    16'd34280: out <= 16'h022F;    16'd34281: out <= 16'hFEA6;    16'd34282: out <= 16'hFC8B;    16'd34283: out <= 16'h03BE;
    16'd34284: out <= 16'hFC25;    16'd34285: out <= 16'hFDF1;    16'd34286: out <= 16'hFE64;    16'd34287: out <= 16'h0213;
    16'd34288: out <= 16'hFDD1;    16'd34289: out <= 16'hFDF0;    16'd34290: out <= 16'hFD85;    16'd34291: out <= 16'hFE1F;
    16'd34292: out <= 16'hFABB;    16'd34293: out <= 16'hFF79;    16'd34294: out <= 16'h0688;    16'd34295: out <= 16'h01A3;
    16'd34296: out <= 16'h036B;    16'd34297: out <= 16'h0096;    16'd34298: out <= 16'h0395;    16'd34299: out <= 16'h03C5;
    16'd34300: out <= 16'h03D5;    16'd34301: out <= 16'h038B;    16'd34302: out <= 16'h0115;    16'd34303: out <= 16'h0531;
    16'd34304: out <= 16'hFCC0;    16'd34305: out <= 16'hFCD9;    16'd34306: out <= 16'h0288;    16'd34307: out <= 16'hFC21;
    16'd34308: out <= 16'hFDB5;    16'd34309: out <= 16'hFBC8;    16'd34310: out <= 16'h0364;    16'd34311: out <= 16'hFDFC;
    16'd34312: out <= 16'hFD7A;    16'd34313: out <= 16'h03E3;    16'd34314: out <= 16'h0410;    16'd34315: out <= 16'hF9A9;
    16'd34316: out <= 16'hF93E;    16'd34317: out <= 16'hFD0C;    16'd34318: out <= 16'h0883;    16'd34319: out <= 16'h0652;
    16'd34320: out <= 16'h05BF;    16'd34321: out <= 16'hFB91;    16'd34322: out <= 16'hFE29;    16'd34323: out <= 16'hFF04;
    16'd34324: out <= 16'h008B;    16'd34325: out <= 16'hFBA5;    16'd34326: out <= 16'hFFE3;    16'd34327: out <= 16'h0857;
    16'd34328: out <= 16'h04CA;    16'd34329: out <= 16'h05D2;    16'd34330: out <= 16'h06B9;    16'd34331: out <= 16'h02BC;
    16'd34332: out <= 16'h0A1C;    16'd34333: out <= 16'hFD41;    16'd34334: out <= 16'hFE2F;    16'd34335: out <= 16'h00BD;
    16'd34336: out <= 16'h02E1;    16'd34337: out <= 16'h0540;    16'd34338: out <= 16'h0850;    16'd34339: out <= 16'h066E;
    16'd34340: out <= 16'h02FB;    16'd34341: out <= 16'h01C5;    16'd34342: out <= 16'h024F;    16'd34343: out <= 16'hFFBC;
    16'd34344: out <= 16'h06D9;    16'd34345: out <= 16'h0371;    16'd34346: out <= 16'h053E;    16'd34347: out <= 16'h05D4;
    16'd34348: out <= 16'h0849;    16'd34349: out <= 16'h06F6;    16'd34350: out <= 16'h0668;    16'd34351: out <= 16'h01D4;
    16'd34352: out <= 16'h01E1;    16'd34353: out <= 16'h028F;    16'd34354: out <= 16'h03BC;    16'd34355: out <= 16'h062F;
    16'd34356: out <= 16'hFC76;    16'd34357: out <= 16'h0273;    16'd34358: out <= 16'h0337;    16'd34359: out <= 16'h06C8;
    16'd34360: out <= 16'h061C;    16'd34361: out <= 16'hFD5B;    16'd34362: out <= 16'h0B99;    16'd34363: out <= 16'h0542;
    16'd34364: out <= 16'h00F6;    16'd34365: out <= 16'h03F6;    16'd34366: out <= 16'h05FF;    16'd34367: out <= 16'h0118;
    16'd34368: out <= 16'h017B;    16'd34369: out <= 16'hFFC0;    16'd34370: out <= 16'h02D4;    16'd34371: out <= 16'h0413;
    16'd34372: out <= 16'h0103;    16'd34373: out <= 16'h0284;    16'd34374: out <= 16'h0763;    16'd34375: out <= 16'h043F;
    16'd34376: out <= 16'h00D1;    16'd34377: out <= 16'hFFB6;    16'd34378: out <= 16'h05D5;    16'd34379: out <= 16'hFACE;
    16'd34380: out <= 16'h0947;    16'd34381: out <= 16'hFE72;    16'd34382: out <= 16'h03D7;    16'd34383: out <= 16'h09E9;
    16'd34384: out <= 16'h01EA;    16'd34385: out <= 16'h0101;    16'd34386: out <= 16'h0236;    16'd34387: out <= 16'h0652;
    16'd34388: out <= 16'h00CB;    16'd34389: out <= 16'h0330;    16'd34390: out <= 16'h0387;    16'd34391: out <= 16'h001F;
    16'd34392: out <= 16'hFEF9;    16'd34393: out <= 16'h02EA;    16'd34394: out <= 16'h032E;    16'd34395: out <= 16'h04CB;
    16'd34396: out <= 16'h06EE;    16'd34397: out <= 16'h0370;    16'd34398: out <= 16'h0369;    16'd34399: out <= 16'h0409;
    16'd34400: out <= 16'h0899;    16'd34401: out <= 16'h045E;    16'd34402: out <= 16'h065E;    16'd34403: out <= 16'h0C3F;
    16'd34404: out <= 16'h02FB;    16'd34405: out <= 16'h0699;    16'd34406: out <= 16'h06DA;    16'd34407: out <= 16'hFD6C;
    16'd34408: out <= 16'h0898;    16'd34409: out <= 16'h02DE;    16'd34410: out <= 16'h0094;    16'd34411: out <= 16'h00E9;
    16'd34412: out <= 16'h0269;    16'd34413: out <= 16'h03AF;    16'd34414: out <= 16'h05F6;    16'd34415: out <= 16'h08A8;
    16'd34416: out <= 16'h0008;    16'd34417: out <= 16'h0664;    16'd34418: out <= 16'h0678;    16'd34419: out <= 16'h0951;
    16'd34420: out <= 16'h01D6;    16'd34421: out <= 16'h0220;    16'd34422: out <= 16'h0616;    16'd34423: out <= 16'h002F;
    16'd34424: out <= 16'h02DF;    16'd34425: out <= 16'h07A2;    16'd34426: out <= 16'h06C5;    16'd34427: out <= 16'h0782;
    16'd34428: out <= 16'h04EB;    16'd34429: out <= 16'h057B;    16'd34430: out <= 16'h06DF;    16'd34431: out <= 16'h0237;
    16'd34432: out <= 16'hFDD8;    16'd34433: out <= 16'h05F9;    16'd34434: out <= 16'hFE9F;    16'd34435: out <= 16'h0598;
    16'd34436: out <= 16'h0488;    16'd34437: out <= 16'h0495;    16'd34438: out <= 16'h017E;    16'd34439: out <= 16'h0223;
    16'd34440: out <= 16'h0781;    16'd34441: out <= 16'h00BF;    16'd34442: out <= 16'h0414;    16'd34443: out <= 16'h0856;
    16'd34444: out <= 16'h0430;    16'd34445: out <= 16'h054A;    16'd34446: out <= 16'h0B46;    16'd34447: out <= 16'hFBDB;
    16'd34448: out <= 16'h008D;    16'd34449: out <= 16'hFF87;    16'd34450: out <= 16'h0815;    16'd34451: out <= 16'h05D5;
    16'd34452: out <= 16'h09AB;    16'd34453: out <= 16'h0A44;    16'd34454: out <= 16'h0075;    16'd34455: out <= 16'h0498;
    16'd34456: out <= 16'h0402;    16'd34457: out <= 16'hFE1B;    16'd34458: out <= 16'h01C2;    16'd34459: out <= 16'h0239;
    16'd34460: out <= 16'h02CE;    16'd34461: out <= 16'h03B7;    16'd34462: out <= 16'h0C6F;    16'd34463: out <= 16'h03CB;
    16'd34464: out <= 16'hFFAA;    16'd34465: out <= 16'h0493;    16'd34466: out <= 16'h084C;    16'd34467: out <= 16'h01A3;
    16'd34468: out <= 16'hFFDA;    16'd34469: out <= 16'h02A7;    16'd34470: out <= 16'hFDB5;    16'd34471: out <= 16'h0775;
    16'd34472: out <= 16'h035B;    16'd34473: out <= 16'h03ED;    16'd34474: out <= 16'h091E;    16'd34475: out <= 16'hFBE1;
    16'd34476: out <= 16'h09D5;    16'd34477: out <= 16'h024B;    16'd34478: out <= 16'h029D;    16'd34479: out <= 16'h04BE;
    16'd34480: out <= 16'h0627;    16'd34481: out <= 16'hFF07;    16'd34482: out <= 16'h0095;    16'd34483: out <= 16'h0772;
    16'd34484: out <= 16'hFE00;    16'd34485: out <= 16'h083C;    16'd34486: out <= 16'h0169;    16'd34487: out <= 16'hFB9C;
    16'd34488: out <= 16'h03C1;    16'd34489: out <= 16'h05AC;    16'd34490: out <= 16'h053A;    16'd34491: out <= 16'h0CBA;
    16'd34492: out <= 16'h013C;    16'd34493: out <= 16'h0055;    16'd34494: out <= 16'h04C4;    16'd34495: out <= 16'h06C8;
    16'd34496: out <= 16'h004F;    16'd34497: out <= 16'h01B6;    16'd34498: out <= 16'h0463;    16'd34499: out <= 16'h033A;
    16'd34500: out <= 16'h02F2;    16'd34501: out <= 16'h04CE;    16'd34502: out <= 16'hFD17;    16'd34503: out <= 16'h05FA;
    16'd34504: out <= 16'hFD41;    16'd34505: out <= 16'h0575;    16'd34506: out <= 16'h0483;    16'd34507: out <= 16'h0125;
    16'd34508: out <= 16'h0486;    16'd34509: out <= 16'h0254;    16'd34510: out <= 16'h07CD;    16'd34511: out <= 16'h03D2;
    16'd34512: out <= 16'h04CB;    16'd34513: out <= 16'hFEF9;    16'd34514: out <= 16'h05FD;    16'd34515: out <= 16'h0AFA;
    16'd34516: out <= 16'h016F;    16'd34517: out <= 16'h004B;    16'd34518: out <= 16'h0099;    16'd34519: out <= 16'h04F5;
    16'd34520: out <= 16'h0152;    16'd34521: out <= 16'h004E;    16'd34522: out <= 16'hFAD5;    16'd34523: out <= 16'h04BB;
    16'd34524: out <= 16'h04DB;    16'd34525: out <= 16'h0067;    16'd34526: out <= 16'h0731;    16'd34527: out <= 16'hFF77;
    16'd34528: out <= 16'h0872;    16'd34529: out <= 16'h0A1A;    16'd34530: out <= 16'h0A64;    16'd34531: out <= 16'h07BA;
    16'd34532: out <= 16'hFB84;    16'd34533: out <= 16'h0006;    16'd34534: out <= 16'hF5EC;    16'd34535: out <= 16'h07C2;
    16'd34536: out <= 16'hFB58;    16'd34537: out <= 16'hFDBC;    16'd34538: out <= 16'h04A5;    16'd34539: out <= 16'hFD93;
    16'd34540: out <= 16'h001D;    16'd34541: out <= 16'h01D1;    16'd34542: out <= 16'h00B9;    16'd34543: out <= 16'h0112;
    16'd34544: out <= 16'h06E1;    16'd34545: out <= 16'h0267;    16'd34546: out <= 16'hFF61;    16'd34547: out <= 16'hFDD4;
    16'd34548: out <= 16'hF904;    16'd34549: out <= 16'h06DC;    16'd34550: out <= 16'h00D1;    16'd34551: out <= 16'hFBFC;
    16'd34552: out <= 16'hFFF4;    16'd34553: out <= 16'h027E;    16'd34554: out <= 16'h01E7;    16'd34555: out <= 16'h026C;
    16'd34556: out <= 16'h0445;    16'd34557: out <= 16'hF6B2;    16'd34558: out <= 16'h04F7;    16'd34559: out <= 16'h01D2;
    16'd34560: out <= 16'hFFE8;    16'd34561: out <= 16'hFD94;    16'd34562: out <= 16'hFFFF;    16'd34563: out <= 16'hFEEC;
    16'd34564: out <= 16'h0849;    16'd34565: out <= 16'h02CD;    16'd34566: out <= 16'h002E;    16'd34567: out <= 16'h0775;
    16'd34568: out <= 16'hFF47;    16'd34569: out <= 16'h0959;    16'd34570: out <= 16'h074E;    16'd34571: out <= 16'hFF76;
    16'd34572: out <= 16'hFC77;    16'd34573: out <= 16'h0114;    16'd34574: out <= 16'hFFEE;    16'd34575: out <= 16'h0274;
    16'd34576: out <= 16'hFD16;    16'd34577: out <= 16'hF80D;    16'd34578: out <= 16'hFAD7;    16'd34579: out <= 16'h0296;
    16'd34580: out <= 16'hFD34;    16'd34581: out <= 16'hFD81;    16'd34582: out <= 16'h01E2;    16'd34583: out <= 16'h0174;
    16'd34584: out <= 16'h0425;    16'd34585: out <= 16'h0784;    16'd34586: out <= 16'h081A;    16'd34587: out <= 16'h0660;
    16'd34588: out <= 16'h01D5;    16'd34589: out <= 16'h0247;    16'd34590: out <= 16'h0398;    16'd34591: out <= 16'h0527;
    16'd34592: out <= 16'h0926;    16'd34593: out <= 16'h051C;    16'd34594: out <= 16'h0833;    16'd34595: out <= 16'hFB9D;
    16'd34596: out <= 16'h060F;    16'd34597: out <= 16'h0A0D;    16'd34598: out <= 16'h06C3;    16'd34599: out <= 16'h0265;
    16'd34600: out <= 16'h0614;    16'd34601: out <= 16'h05F4;    16'd34602: out <= 16'h0288;    16'd34603: out <= 16'h0A87;
    16'd34604: out <= 16'h06A1;    16'd34605: out <= 16'h0904;    16'd34606: out <= 16'hFF9D;    16'd34607: out <= 16'h0477;
    16'd34608: out <= 16'h02E1;    16'd34609: out <= 16'h02A9;    16'd34610: out <= 16'h0975;    16'd34611: out <= 16'hFE7C;
    16'd34612: out <= 16'h0373;    16'd34613: out <= 16'hFA4A;    16'd34614: out <= 16'h01F7;    16'd34615: out <= 16'h06CD;
    16'd34616: out <= 16'h041E;    16'd34617: out <= 16'h0627;    16'd34618: out <= 16'h0A84;    16'd34619: out <= 16'h0C0A;
    16'd34620: out <= 16'h05BF;    16'd34621: out <= 16'h0271;    16'd34622: out <= 16'h09EB;    16'd34623: out <= 16'h0653;
    16'd34624: out <= 16'h0194;    16'd34625: out <= 16'hFEF6;    16'd34626: out <= 16'h03D4;    16'd34627: out <= 16'h0377;
    16'd34628: out <= 16'h06DA;    16'd34629: out <= 16'h00C3;    16'd34630: out <= 16'h03A0;    16'd34631: out <= 16'h00FC;
    16'd34632: out <= 16'h03C0;    16'd34633: out <= 16'h06F2;    16'd34634: out <= 16'hFD63;    16'd34635: out <= 16'h0286;
    16'd34636: out <= 16'h049F;    16'd34637: out <= 16'hFBA2;    16'd34638: out <= 16'h00AB;    16'd34639: out <= 16'h0951;
    16'd34640: out <= 16'h046B;    16'd34641: out <= 16'h003E;    16'd34642: out <= 16'h0185;    16'd34643: out <= 16'h076D;
    16'd34644: out <= 16'h0463;    16'd34645: out <= 16'h02F0;    16'd34646: out <= 16'h08A3;    16'd34647: out <= 16'h07AA;
    16'd34648: out <= 16'h0CAA;    16'd34649: out <= 16'h01D6;    16'd34650: out <= 16'h05A5;    16'd34651: out <= 16'h02B4;
    16'd34652: out <= 16'h0600;    16'd34653: out <= 16'h0992;    16'd34654: out <= 16'h009C;    16'd34655: out <= 16'h02ED;
    16'd34656: out <= 16'h0289;    16'd34657: out <= 16'h069F;    16'd34658: out <= 16'h02F8;    16'd34659: out <= 16'hFFE6;
    16'd34660: out <= 16'h0BBC;    16'd34661: out <= 16'h00B9;    16'd34662: out <= 16'h00C9;    16'd34663: out <= 16'h03C0;
    16'd34664: out <= 16'hFE61;    16'd34665: out <= 16'hFF60;    16'd34666: out <= 16'hFB0A;    16'd34667: out <= 16'h02FC;
    16'd34668: out <= 16'h05B9;    16'd34669: out <= 16'hFD94;    16'd34670: out <= 16'hFF4F;    16'd34671: out <= 16'h0440;
    16'd34672: out <= 16'hFE8C;    16'd34673: out <= 16'h0449;    16'd34674: out <= 16'h0495;    16'd34675: out <= 16'hFDB7;
    16'd34676: out <= 16'h04DA;    16'd34677: out <= 16'h081F;    16'd34678: out <= 16'h0059;    16'd34679: out <= 16'h00FE;
    16'd34680: out <= 16'h066F;    16'd34681: out <= 16'h05E0;    16'd34682: out <= 16'h0889;    16'd34683: out <= 16'h0561;
    16'd34684: out <= 16'h00E3;    16'd34685: out <= 16'h0669;    16'd34686: out <= 16'h060A;    16'd34687: out <= 16'h02CA;
    16'd34688: out <= 16'h0ABE;    16'd34689: out <= 16'h05CC;    16'd34690: out <= 16'h02AC;    16'd34691: out <= 16'h052D;
    16'd34692: out <= 16'hFEDF;    16'd34693: out <= 16'h01AA;    16'd34694: out <= 16'h0ABF;    16'd34695: out <= 16'h03C1;
    16'd34696: out <= 16'hFFC4;    16'd34697: out <= 16'h11E5;    16'd34698: out <= 16'h0033;    16'd34699: out <= 16'h04F2;
    16'd34700: out <= 16'h0006;    16'd34701: out <= 16'h08FC;    16'd34702: out <= 16'hFC82;    16'd34703: out <= 16'h0777;
    16'd34704: out <= 16'h0656;    16'd34705: out <= 16'h03A3;    16'd34706: out <= 16'h092A;    16'd34707: out <= 16'h02B8;
    16'd34708: out <= 16'h0620;    16'd34709: out <= 16'h00FC;    16'd34710: out <= 16'h023E;    16'd34711: out <= 16'h0639;
    16'd34712: out <= 16'h0226;    16'd34713: out <= 16'h0443;    16'd34714: out <= 16'h067E;    16'd34715: out <= 16'h06C4;
    16'd34716: out <= 16'h02B9;    16'd34717: out <= 16'h078A;    16'd34718: out <= 16'h05FA;    16'd34719: out <= 16'h097F;
    16'd34720: out <= 16'h05FF;    16'd34721: out <= 16'hFE57;    16'd34722: out <= 16'h0471;    16'd34723: out <= 16'hFD77;
    16'd34724: out <= 16'h0F55;    16'd34725: out <= 16'h05EE;    16'd34726: out <= 16'hF715;    16'd34727: out <= 16'h00F8;
    16'd34728: out <= 16'h015B;    16'd34729: out <= 16'h002E;    16'd34730: out <= 16'h015F;    16'd34731: out <= 16'h019F;
    16'd34732: out <= 16'hF8EA;    16'd34733: out <= 16'h0478;    16'd34734: out <= 16'h00DD;    16'd34735: out <= 16'hFCDD;
    16'd34736: out <= 16'hFFDE;    16'd34737: out <= 16'h0723;    16'd34738: out <= 16'h030A;    16'd34739: out <= 16'hFD40;
    16'd34740: out <= 16'h08C4;    16'd34741: out <= 16'h04E6;    16'd34742: out <= 16'h05FA;    16'd34743: out <= 16'h011D;
    16'd34744: out <= 16'h0667;    16'd34745: out <= 16'hFC9C;    16'd34746: out <= 16'h083E;    16'd34747: out <= 16'h0158;
    16'd34748: out <= 16'h02DC;    16'd34749: out <= 16'h00B3;    16'd34750: out <= 16'h07A0;    16'd34751: out <= 16'h0B5D;
    16'd34752: out <= 16'h0776;    16'd34753: out <= 16'h024E;    16'd34754: out <= 16'h03F9;    16'd34755: out <= 16'h039E;
    16'd34756: out <= 16'h0B0D;    16'd34757: out <= 16'hFC9A;    16'd34758: out <= 16'h049F;    16'd34759: out <= 16'h05E1;
    16'd34760: out <= 16'h025E;    16'd34761: out <= 16'hFD70;    16'd34762: out <= 16'h0062;    16'd34763: out <= 16'h031E;
    16'd34764: out <= 16'h0403;    16'd34765: out <= 16'h0271;    16'd34766: out <= 16'h00B4;    16'd34767: out <= 16'h044F;
    16'd34768: out <= 16'h0103;    16'd34769: out <= 16'h00FB;    16'd34770: out <= 16'h060B;    16'd34771: out <= 16'h00E7;
    16'd34772: out <= 16'h0530;    16'd34773: out <= 16'h03D3;    16'd34774: out <= 16'h07BF;    16'd34775: out <= 16'hFF46;
    16'd34776: out <= 16'h03EA;    16'd34777: out <= 16'hF8EA;    16'd34778: out <= 16'h00EC;    16'd34779: out <= 16'h0A3F;
    16'd34780: out <= 16'hFE65;    16'd34781: out <= 16'h0431;    16'd34782: out <= 16'h07B2;    16'd34783: out <= 16'h05FA;
    16'd34784: out <= 16'h09F7;    16'd34785: out <= 16'h031E;    16'd34786: out <= 16'hFE52;    16'd34787: out <= 16'h043F;
    16'd34788: out <= 16'h0554;    16'd34789: out <= 16'hFB5F;    16'd34790: out <= 16'hFC0E;    16'd34791: out <= 16'h04E9;
    16'd34792: out <= 16'hFC98;    16'd34793: out <= 16'h038F;    16'd34794: out <= 16'h039D;    16'd34795: out <= 16'hFDE4;
    16'd34796: out <= 16'hFF34;    16'd34797: out <= 16'h0131;    16'd34798: out <= 16'hFB95;    16'd34799: out <= 16'h0396;
    16'd34800: out <= 16'h039B;    16'd34801: out <= 16'hFF52;    16'd34802: out <= 16'hFFDF;    16'd34803: out <= 16'h02BF;
    16'd34804: out <= 16'hF7B4;    16'd34805: out <= 16'h01D9;    16'd34806: out <= 16'hFE7C;    16'd34807: out <= 16'h031F;
    16'd34808: out <= 16'hFD7E;    16'd34809: out <= 16'h0000;    16'd34810: out <= 16'h00B7;    16'd34811: out <= 16'h03FA;
    16'd34812: out <= 16'hFF12;    16'd34813: out <= 16'h0257;    16'd34814: out <= 16'h0360;    16'd34815: out <= 16'hFEB0;
    16'd34816: out <= 16'h03F4;    16'd34817: out <= 16'hFE9F;    16'd34818: out <= 16'h0117;    16'd34819: out <= 16'hFD4C;
    16'd34820: out <= 16'h0126;    16'd34821: out <= 16'h07E6;    16'd34822: out <= 16'hFFBF;    16'd34823: out <= 16'h0434;
    16'd34824: out <= 16'hFE56;    16'd34825: out <= 16'hFEF7;    16'd34826: out <= 16'hF6FD;    16'd34827: out <= 16'hFBEF;
    16'd34828: out <= 16'h0150;    16'd34829: out <= 16'hFACA;    16'd34830: out <= 16'h065C;    16'd34831: out <= 16'hFD9D;
    16'd34832: out <= 16'h00A2;    16'd34833: out <= 16'h014E;    16'd34834: out <= 16'h00BB;    16'd34835: out <= 16'hFD0E;
    16'd34836: out <= 16'hFC9D;    16'd34837: out <= 16'hFD6D;    16'd34838: out <= 16'h0158;    16'd34839: out <= 16'h0137;
    16'd34840: out <= 16'h02E3;    16'd34841: out <= 16'h05F2;    16'd34842: out <= 16'h0023;    16'd34843: out <= 16'h0088;
    16'd34844: out <= 16'hFD44;    16'd34845: out <= 16'h02FE;    16'd34846: out <= 16'h02EA;    16'd34847: out <= 16'h055F;
    16'd34848: out <= 16'hFEC1;    16'd34849: out <= 16'h03E4;    16'd34850: out <= 16'h00EA;    16'd34851: out <= 16'h0810;
    16'd34852: out <= 16'h0445;    16'd34853: out <= 16'h0176;    16'd34854: out <= 16'h09C9;    16'd34855: out <= 16'h0488;
    16'd34856: out <= 16'h0412;    16'd34857: out <= 16'h03ED;    16'd34858: out <= 16'h053A;    16'd34859: out <= 16'hFCCC;
    16'd34860: out <= 16'h01D3;    16'd34861: out <= 16'h06A0;    16'd34862: out <= 16'h00A1;    16'd34863: out <= 16'hFED3;
    16'd34864: out <= 16'hFAF8;    16'd34865: out <= 16'h0056;    16'd34866: out <= 16'h03C4;    16'd34867: out <= 16'h0180;
    16'd34868: out <= 16'h032A;    16'd34869: out <= 16'h0763;    16'd34870: out <= 16'h072E;    16'd34871: out <= 16'h03F8;
    16'd34872: out <= 16'h0655;    16'd34873: out <= 16'h0380;    16'd34874: out <= 16'h0516;    16'd34875: out <= 16'h077C;
    16'd34876: out <= 16'h0458;    16'd34877: out <= 16'h0644;    16'd34878: out <= 16'h08FB;    16'd34879: out <= 16'h03BB;
    16'd34880: out <= 16'h0152;    16'd34881: out <= 16'h0584;    16'd34882: out <= 16'h021F;    16'd34883: out <= 16'h0EE7;
    16'd34884: out <= 16'h0563;    16'd34885: out <= 16'h042C;    16'd34886: out <= 16'h0488;    16'd34887: out <= 16'h039F;
    16'd34888: out <= 16'h09CA;    16'd34889: out <= 16'h04F0;    16'd34890: out <= 16'h062D;    16'd34891: out <= 16'h0293;
    16'd34892: out <= 16'h042C;    16'd34893: out <= 16'h0754;    16'd34894: out <= 16'hFBEE;    16'd34895: out <= 16'h0636;
    16'd34896: out <= 16'h02C6;    16'd34897: out <= 16'h036D;    16'd34898: out <= 16'h068B;    16'd34899: out <= 16'h06AD;
    16'd34900: out <= 16'hFE04;    16'd34901: out <= 16'h029F;    16'd34902: out <= 16'h01AF;    16'd34903: out <= 16'h09A2;
    16'd34904: out <= 16'h08DB;    16'd34905: out <= 16'h0182;    16'd34906: out <= 16'h026E;    16'd34907: out <= 16'h0718;
    16'd34908: out <= 16'h0693;    16'd34909: out <= 16'hFFD4;    16'd34910: out <= 16'h0222;    16'd34911: out <= 16'h05BF;
    16'd34912: out <= 16'h027F;    16'd34913: out <= 16'h05E0;    16'd34914: out <= 16'h06A6;    16'd34915: out <= 16'hFD8E;
    16'd34916: out <= 16'hFFD5;    16'd34917: out <= 16'h000C;    16'd34918: out <= 16'h0867;    16'd34919: out <= 16'h098A;
    16'd34920: out <= 16'h0546;    16'd34921: out <= 16'h0336;    16'd34922: out <= 16'h057B;    16'd34923: out <= 16'h0574;
    16'd34924: out <= 16'h04D9;    16'd34925: out <= 16'h044D;    16'd34926: out <= 16'h0799;    16'd34927: out <= 16'h0303;
    16'd34928: out <= 16'h044F;    16'd34929: out <= 16'h0350;    16'd34930: out <= 16'h0162;    16'd34931: out <= 16'h0254;
    16'd34932: out <= 16'h04C6;    16'd34933: out <= 16'h050D;    16'd34934: out <= 16'h02A8;    16'd34935: out <= 16'h08F3;
    16'd34936: out <= 16'h0236;    16'd34937: out <= 16'h072F;    16'd34938: out <= 16'h03FE;    16'd34939: out <= 16'h0C0A;
    16'd34940: out <= 16'hFF19;    16'd34941: out <= 16'h0CD6;    16'd34942: out <= 16'hFEDB;    16'd34943: out <= 16'h02BC;
    16'd34944: out <= 16'h033C;    16'd34945: out <= 16'h0690;    16'd34946: out <= 16'h0394;    16'd34947: out <= 16'h039B;
    16'd34948: out <= 16'hFE09;    16'd34949: out <= 16'h0475;    16'd34950: out <= 16'h097A;    16'd34951: out <= 16'h03A6;
    16'd34952: out <= 16'h0D18;    16'd34953: out <= 16'h03FD;    16'd34954: out <= 16'h069D;    16'd34955: out <= 16'h08C8;
    16'd34956: out <= 16'h0213;    16'd34957: out <= 16'h0379;    16'd34958: out <= 16'h0968;    16'd34959: out <= 16'h069A;
    16'd34960: out <= 16'h03EA;    16'd34961: out <= 16'h071D;    16'd34962: out <= 16'h0395;    16'd34963: out <= 16'h0558;
    16'd34964: out <= 16'h05BF;    16'd34965: out <= 16'h071B;    16'd34966: out <= 16'h0627;    16'd34967: out <= 16'h05ED;
    16'd34968: out <= 16'h0364;    16'd34969: out <= 16'h0030;    16'd34970: out <= 16'hFCEF;    16'd34971: out <= 16'h0254;
    16'd34972: out <= 16'h0789;    16'd34973: out <= 16'h0375;    16'd34974: out <= 16'hFD62;    16'd34975: out <= 16'hFF50;
    16'd34976: out <= 16'h01E5;    16'd34977: out <= 16'h0386;    16'd34978: out <= 16'h034D;    16'd34979: out <= 16'hFE3D;
    16'd34980: out <= 16'hFEAC;    16'd34981: out <= 16'h05FA;    16'd34982: out <= 16'hFEBB;    16'd34983: out <= 16'h0769;
    16'd34984: out <= 16'h0630;    16'd34985: out <= 16'h0722;    16'd34986: out <= 16'h0393;    16'd34987: out <= 16'h0741;
    16'd34988: out <= 16'h0405;    16'd34989: out <= 16'hFF68;    16'd34990: out <= 16'h073A;    16'd34991: out <= 16'h00DA;
    16'd34992: out <= 16'hFAA3;    16'd34993: out <= 16'h06EB;    16'd34994: out <= 16'h0626;    16'd34995: out <= 16'h0465;
    16'd34996: out <= 16'h0853;    16'd34997: out <= 16'h0235;    16'd34998: out <= 16'hFFE5;    16'd34999: out <= 16'hFEB8;
    16'd35000: out <= 16'h0329;    16'd35001: out <= 16'h04D7;    16'd35002: out <= 16'hFF0F;    16'd35003: out <= 16'hFC0D;
    16'd35004: out <= 16'h030D;    16'd35005: out <= 16'h0635;    16'd35006: out <= 16'h00A2;    16'd35007: out <= 16'h046E;
    16'd35008: out <= 16'h03CE;    16'd35009: out <= 16'h03C5;    16'd35010: out <= 16'h03BC;    16'd35011: out <= 16'h0239;
    16'd35012: out <= 16'h02FA;    16'd35013: out <= 16'h05B2;    16'd35014: out <= 16'hFFEF;    16'd35015: out <= 16'h0282;
    16'd35016: out <= 16'h0575;    16'd35017: out <= 16'h02C5;    16'd35018: out <= 16'h0836;    16'd35019: out <= 16'hFFCA;
    16'd35020: out <= 16'hFF38;    16'd35021: out <= 16'h024A;    16'd35022: out <= 16'hFB8D;    16'd35023: out <= 16'h025C;
    16'd35024: out <= 16'h00F0;    16'd35025: out <= 16'h0645;    16'd35026: out <= 16'h0C43;    16'd35027: out <= 16'h039D;
    16'd35028: out <= 16'h0301;    16'd35029: out <= 16'h05FA;    16'd35030: out <= 16'h0655;    16'd35031: out <= 16'h032D;
    16'd35032: out <= 16'hFC09;    16'd35033: out <= 16'h0245;    16'd35034: out <= 16'h02D2;    16'd35035: out <= 16'hFFBF;
    16'd35036: out <= 16'h0171;    16'd35037: out <= 16'hFD5E;    16'd35038: out <= 16'h043D;    16'd35039: out <= 16'h04D4;
    16'd35040: out <= 16'h0707;    16'd35041: out <= 16'hFD40;    16'd35042: out <= 16'h0424;    16'd35043: out <= 16'h00F8;
    16'd35044: out <= 16'h0B54;    16'd35045: out <= 16'h07B0;    16'd35046: out <= 16'h03A7;    16'd35047: out <= 16'h0411;
    16'd35048: out <= 16'h0478;    16'd35049: out <= 16'hFA71;    16'd35050: out <= 16'hFB2B;    16'd35051: out <= 16'hF903;
    16'd35052: out <= 16'h0040;    16'd35053: out <= 16'h01F1;    16'd35054: out <= 16'hF9CA;    16'd35055: out <= 16'h06C4;
    16'd35056: out <= 16'h062C;    16'd35057: out <= 16'hFB3C;    16'd35058: out <= 16'h09A6;    16'd35059: out <= 16'h0041;
    16'd35060: out <= 16'h0100;    16'd35061: out <= 16'hFD33;    16'd35062: out <= 16'h031B;    16'd35063: out <= 16'hFD1B;
    16'd35064: out <= 16'hFD8E;    16'd35065: out <= 16'hFC44;    16'd35066: out <= 16'h01C3;    16'd35067: out <= 16'h0376;
    16'd35068: out <= 16'hF99F;    16'd35069: out <= 16'h047E;    16'd35070: out <= 16'h049E;    16'd35071: out <= 16'hFE0F;
    16'd35072: out <= 16'hFEBE;    16'd35073: out <= 16'hFD5A;    16'd35074: out <= 16'h0631;    16'd35075: out <= 16'hFCD8;
    16'd35076: out <= 16'hFF71;    16'd35077: out <= 16'h00AF;    16'd35078: out <= 16'h0637;    16'd35079: out <= 16'hFFCA;
    16'd35080: out <= 16'hFE60;    16'd35081: out <= 16'h02F8;    16'd35082: out <= 16'h050D;    16'd35083: out <= 16'h01DE;
    16'd35084: out <= 16'h0483;    16'd35085: out <= 16'h06B6;    16'd35086: out <= 16'hFC17;    16'd35087: out <= 16'hFF2E;
    16'd35088: out <= 16'hFF8C;    16'd35089: out <= 16'h015D;    16'd35090: out <= 16'hF7F3;    16'd35091: out <= 16'h022B;
    16'd35092: out <= 16'hFEA2;    16'd35093: out <= 16'h0004;    16'd35094: out <= 16'hFF7B;    16'd35095: out <= 16'hFFB9;
    16'd35096: out <= 16'h07CD;    16'd35097: out <= 16'h009F;    16'd35098: out <= 16'hFE69;    16'd35099: out <= 16'h0310;
    16'd35100: out <= 16'h00F2;    16'd35101: out <= 16'h015C;    16'd35102: out <= 16'h03C3;    16'd35103: out <= 16'h08E3;
    16'd35104: out <= 16'h067F;    16'd35105: out <= 16'h029C;    16'd35106: out <= 16'h051B;    16'd35107: out <= 16'h02B9;
    16'd35108: out <= 16'h009B;    16'd35109: out <= 16'h04CE;    16'd35110: out <= 16'h04AB;    16'd35111: out <= 16'h04AC;
    16'd35112: out <= 16'h0785;    16'd35113: out <= 16'h016D;    16'd35114: out <= 16'hFBC7;    16'd35115: out <= 16'h0907;
    16'd35116: out <= 16'h0388;    16'd35117: out <= 16'h01D9;    16'd35118: out <= 16'h0336;    16'd35119: out <= 16'h04AB;
    16'd35120: out <= 16'hFD5D;    16'd35121: out <= 16'h024B;    16'd35122: out <= 16'h0386;    16'd35123: out <= 16'h0799;
    16'd35124: out <= 16'hFEC8;    16'd35125: out <= 16'hFF3E;    16'd35126: out <= 16'h08F5;    16'd35127: out <= 16'hFD69;
    16'd35128: out <= 16'h029B;    16'd35129: out <= 16'h0C26;    16'd35130: out <= 16'h0245;    16'd35131: out <= 16'hFDA3;
    16'd35132: out <= 16'hFF61;    16'd35133: out <= 16'h0218;    16'd35134: out <= 16'h047C;    16'd35135: out <= 16'h0026;
    16'd35136: out <= 16'h05DF;    16'd35137: out <= 16'h0D70;    16'd35138: out <= 16'h00CD;    16'd35139: out <= 16'h0929;
    16'd35140: out <= 16'hFFD2;    16'd35141: out <= 16'h0A49;    16'd35142: out <= 16'h0628;    16'd35143: out <= 16'h0AC5;
    16'd35144: out <= 16'hFF37;    16'd35145: out <= 16'h02E8;    16'd35146: out <= 16'h0C9F;    16'd35147: out <= 16'hFF0F;
    16'd35148: out <= 16'h040F;    16'd35149: out <= 16'h0470;    16'd35150: out <= 16'h0B5B;    16'd35151: out <= 16'h0986;
    16'd35152: out <= 16'h02DE;    16'd35153: out <= 16'h0522;    16'd35154: out <= 16'h087E;    16'd35155: out <= 16'h0B59;
    16'd35156: out <= 16'h076E;    16'd35157: out <= 16'hFFA7;    16'd35158: out <= 16'h058B;    16'd35159: out <= 16'h09C9;
    16'd35160: out <= 16'h046E;    16'd35161: out <= 16'hFDB2;    16'd35162: out <= 16'h0247;    16'd35163: out <= 16'h055D;
    16'd35164: out <= 16'h00F5;    16'd35165: out <= 16'h022F;    16'd35166: out <= 16'h0346;    16'd35167: out <= 16'h0671;
    16'd35168: out <= 16'h06AF;    16'd35169: out <= 16'h044D;    16'd35170: out <= 16'h0A20;    16'd35171: out <= 16'h028B;
    16'd35172: out <= 16'h05FA;    16'd35173: out <= 16'h0327;    16'd35174: out <= 16'hFE7A;    16'd35175: out <= 16'h0722;
    16'd35176: out <= 16'h08CF;    16'd35177: out <= 16'h020F;    16'd35178: out <= 16'h0410;    16'd35179: out <= 16'h05CD;
    16'd35180: out <= 16'h04BD;    16'd35181: out <= 16'h0D27;    16'd35182: out <= 16'h05C9;    16'd35183: out <= 16'h08B3;
    16'd35184: out <= 16'h0152;    16'd35185: out <= 16'h028B;    16'd35186: out <= 16'hFFC7;    16'd35187: out <= 16'h01E3;
    16'd35188: out <= 16'h01D9;    16'd35189: out <= 16'h05B4;    16'd35190: out <= 16'h0B2F;    16'd35191: out <= 16'h080E;
    16'd35192: out <= 16'hFE1B;    16'd35193: out <= 16'h0987;    16'd35194: out <= 16'h060A;    16'd35195: out <= 16'h03C0;
    16'd35196: out <= 16'h07F1;    16'd35197: out <= 16'h060A;    16'd35198: out <= 16'h0183;    16'd35199: out <= 16'h079C;
    16'd35200: out <= 16'h0220;    16'd35201: out <= 16'h0234;    16'd35202: out <= 16'h0261;    16'd35203: out <= 16'h0757;
    16'd35204: out <= 16'hFE01;    16'd35205: out <= 16'hFF95;    16'd35206: out <= 16'h0528;    16'd35207: out <= 16'h05CF;
    16'd35208: out <= 16'h09A4;    16'd35209: out <= 16'h0219;    16'd35210: out <= 16'h0CEA;    16'd35211: out <= 16'h0747;
    16'd35212: out <= 16'h0783;    16'd35213: out <= 16'h0053;    16'd35214: out <= 16'h0204;    16'd35215: out <= 16'h0B2C;
    16'd35216: out <= 16'h01CB;    16'd35217: out <= 16'h0015;    16'd35218: out <= 16'hFD90;    16'd35219: out <= 16'h054E;
    16'd35220: out <= 16'h07BE;    16'd35221: out <= 16'h0A08;    16'd35222: out <= 16'h05FB;    16'd35223: out <= 16'h05A5;
    16'd35224: out <= 16'h0521;    16'd35225: out <= 16'h00CF;    16'd35226: out <= 16'h006C;    16'd35227: out <= 16'h0364;
    16'd35228: out <= 16'h06B8;    16'd35229: out <= 16'h070C;    16'd35230: out <= 16'h0376;    16'd35231: out <= 16'h0596;
    16'd35232: out <= 16'h005E;    16'd35233: out <= 16'h0446;    16'd35234: out <= 16'h09DD;    16'd35235: out <= 16'h0799;
    16'd35236: out <= 16'h0391;    16'd35237: out <= 16'h02DF;    16'd35238: out <= 16'h039B;    16'd35239: out <= 16'h04BE;
    16'd35240: out <= 16'h01DF;    16'd35241: out <= 16'h0341;    16'd35242: out <= 16'h04C4;    16'd35243: out <= 16'h00A1;
    16'd35244: out <= 16'h02A2;    16'd35245: out <= 16'h055F;    16'd35246: out <= 16'hFE81;    16'd35247: out <= 16'hFF73;
    16'd35248: out <= 16'h00A3;    16'd35249: out <= 16'h03FE;    16'd35250: out <= 16'h0446;    16'd35251: out <= 16'h0407;
    16'd35252: out <= 16'h064B;    16'd35253: out <= 16'h03D5;    16'd35254: out <= 16'h02F8;    16'd35255: out <= 16'h0101;
    16'd35256: out <= 16'hFFDE;    16'd35257: out <= 16'hFD2A;    16'd35258: out <= 16'h0491;    16'd35259: out <= 16'h0361;
    16'd35260: out <= 16'h03DF;    16'd35261: out <= 16'h00EF;    16'd35262: out <= 16'hFF42;    16'd35263: out <= 16'h026D;
    16'd35264: out <= 16'h01E4;    16'd35265: out <= 16'h032A;    16'd35266: out <= 16'h0443;    16'd35267: out <= 16'h0307;
    16'd35268: out <= 16'h066F;    16'd35269: out <= 16'h0333;    16'd35270: out <= 16'hFC71;    16'd35271: out <= 16'hFC83;
    16'd35272: out <= 16'h04F8;    16'd35273: out <= 16'h0572;    16'd35274: out <= 16'h04BA;    16'd35275: out <= 16'h01F1;
    16'd35276: out <= 16'h0626;    16'd35277: out <= 16'h04C6;    16'd35278: out <= 16'hFB98;    16'd35279: out <= 16'hFDC7;
    16'd35280: out <= 16'h0436;    16'd35281: out <= 16'h07B2;    16'd35282: out <= 16'h02C3;    16'd35283: out <= 16'h05D1;
    16'd35284: out <= 16'h01F7;    16'd35285: out <= 16'hFE0F;    16'd35286: out <= 16'hFBF7;    16'd35287: out <= 16'h019F;
    16'd35288: out <= 16'hFE2D;    16'd35289: out <= 16'hFEE5;    16'd35290: out <= 16'hFE54;    16'd35291: out <= 16'h035E;
    16'd35292: out <= 16'hFDBF;    16'd35293: out <= 16'h03E9;    16'd35294: out <= 16'h0D13;    16'd35295: out <= 16'h04A3;
    16'd35296: out <= 16'h04FC;    16'd35297: out <= 16'hFF2D;    16'd35298: out <= 16'h033A;    16'd35299: out <= 16'h015C;
    16'd35300: out <= 16'h0530;    16'd35301: out <= 16'h0731;    16'd35302: out <= 16'h0455;    16'd35303: out <= 16'hFE89;
    16'd35304: out <= 16'hF7F3;    16'd35305: out <= 16'h00F3;    16'd35306: out <= 16'hFF2E;    16'd35307: out <= 16'h017A;
    16'd35308: out <= 16'hF85A;    16'd35309: out <= 16'hFF0C;    16'd35310: out <= 16'hFB83;    16'd35311: out <= 16'h07C2;
    16'd35312: out <= 16'hFE94;    16'd35313: out <= 16'hF9F1;    16'd35314: out <= 16'h0405;    16'd35315: out <= 16'h003E;
    16'd35316: out <= 16'h071A;    16'd35317: out <= 16'hFEDC;    16'd35318: out <= 16'hFD91;    16'd35319: out <= 16'hF958;
    16'd35320: out <= 16'h000E;    16'd35321: out <= 16'hFE1A;    16'd35322: out <= 16'hFA11;    16'd35323: out <= 16'hFD25;
    16'd35324: out <= 16'hFD24;    16'd35325: out <= 16'h0386;    16'd35326: out <= 16'hFFC8;    16'd35327: out <= 16'h0036;
    16'd35328: out <= 16'h06DD;    16'd35329: out <= 16'hFD58;    16'd35330: out <= 16'hFE76;    16'd35331: out <= 16'h0057;
    16'd35332: out <= 16'hFBEC;    16'd35333: out <= 16'hFB9C;    16'd35334: out <= 16'hFE64;    16'd35335: out <= 16'h02F1;
    16'd35336: out <= 16'hFFD4;    16'd35337: out <= 16'h03DF;    16'd35338: out <= 16'h0314;    16'd35339: out <= 16'h0477;
    16'd35340: out <= 16'h0824;    16'd35341: out <= 16'h0291;    16'd35342: out <= 16'hFC58;    16'd35343: out <= 16'hF681;
    16'd35344: out <= 16'hFE6D;    16'd35345: out <= 16'hFD29;    16'd35346: out <= 16'h01A6;    16'd35347: out <= 16'h0575;
    16'd35348: out <= 16'h02BE;    16'd35349: out <= 16'h04E7;    16'd35350: out <= 16'hF738;    16'd35351: out <= 16'h0189;
    16'd35352: out <= 16'h04F4;    16'd35353: out <= 16'h07BA;    16'd35354: out <= 16'h0963;    16'd35355: out <= 16'h0135;
    16'd35356: out <= 16'h03D0;    16'd35357: out <= 16'h02F7;    16'd35358: out <= 16'h07AE;    16'd35359: out <= 16'hFF23;
    16'd35360: out <= 16'h04A3;    16'd35361: out <= 16'h0420;    16'd35362: out <= 16'h0432;    16'd35363: out <= 16'h0735;
    16'd35364: out <= 16'h02C6;    16'd35365: out <= 16'h01A7;    16'd35366: out <= 16'h0123;    16'd35367: out <= 16'hFFBD;
    16'd35368: out <= 16'h066E;    16'd35369: out <= 16'h02F5;    16'd35370: out <= 16'h0A14;    16'd35371: out <= 16'h01B5;
    16'd35372: out <= 16'h0008;    16'd35373: out <= 16'h0BCD;    16'd35374: out <= 16'h0238;    16'd35375: out <= 16'h0347;
    16'd35376: out <= 16'h0BC7;    16'd35377: out <= 16'h0120;    16'd35378: out <= 16'h054C;    16'd35379: out <= 16'h074B;
    16'd35380: out <= 16'h09ED;    16'd35381: out <= 16'h0E44;    16'd35382: out <= 16'h02FD;    16'd35383: out <= 16'h07FD;
    16'd35384: out <= 16'h041F;    16'd35385: out <= 16'h06D3;    16'd35386: out <= 16'h0664;    16'd35387: out <= 16'h0294;
    16'd35388: out <= 16'h07EC;    16'd35389: out <= 16'h0807;    16'd35390: out <= 16'h081A;    16'd35391: out <= 16'h00F6;
    16'd35392: out <= 16'h0686;    16'd35393: out <= 16'hFEA8;    16'd35394: out <= 16'h0649;    16'd35395: out <= 16'hFA4C;
    16'd35396: out <= 16'h0106;    16'd35397: out <= 16'h027C;    16'd35398: out <= 16'hFD90;    16'd35399: out <= 16'h01ED;
    16'd35400: out <= 16'h003F;    16'd35401: out <= 16'h071C;    16'd35402: out <= 16'h02C7;    16'd35403: out <= 16'h07FF;
    16'd35404: out <= 16'hFFB6;    16'd35405: out <= 16'h09EA;    16'd35406: out <= 16'h04BD;    16'd35407: out <= 16'h0349;
    16'd35408: out <= 16'h0012;    16'd35409: out <= 16'hFD3C;    16'd35410: out <= 16'hFDFA;    16'd35411: out <= 16'h003A;
    16'd35412: out <= 16'h062E;    16'd35413: out <= 16'h0348;    16'd35414: out <= 16'h0A1B;    16'd35415: out <= 16'h025E;
    16'd35416: out <= 16'h01AE;    16'd35417: out <= 16'h0384;    16'd35418: out <= 16'h01BF;    16'd35419: out <= 16'h04BB;
    16'd35420: out <= 16'hFFE7;    16'd35421: out <= 16'h00C1;    16'd35422: out <= 16'h0302;    16'd35423: out <= 16'h0555;
    16'd35424: out <= 16'h062A;    16'd35425: out <= 16'h07A9;    16'd35426: out <= 16'h065E;    16'd35427: out <= 16'h01B4;
    16'd35428: out <= 16'h08A4;    16'd35429: out <= 16'h0344;    16'd35430: out <= 16'hFF00;    16'd35431: out <= 16'hFFAF;
    16'd35432: out <= 16'h058E;    16'd35433: out <= 16'h0B2B;    16'd35434: out <= 16'h07EF;    16'd35435: out <= 16'h00B8;
    16'd35436: out <= 16'h0404;    16'd35437: out <= 16'hFD8A;    16'd35438: out <= 16'h051B;    16'd35439: out <= 16'h0026;
    16'd35440: out <= 16'hFC95;    16'd35441: out <= 16'hFCC6;    16'd35442: out <= 16'h025C;    16'd35443: out <= 16'hFDE2;
    16'd35444: out <= 16'h031E;    16'd35445: out <= 16'h0360;    16'd35446: out <= 16'hFF46;    16'd35447: out <= 16'h06CA;
    16'd35448: out <= 16'h022F;    16'd35449: out <= 16'h08A9;    16'd35450: out <= 16'h0215;    16'd35451: out <= 16'h0210;
    16'd35452: out <= 16'h0F6B;    16'd35453: out <= 16'h0205;    16'd35454: out <= 16'h0743;    16'd35455: out <= 16'h0326;
    16'd35456: out <= 16'h0424;    16'd35457: out <= 16'hFEFA;    16'd35458: out <= 16'h0547;    16'd35459: out <= 16'h00A1;
    16'd35460: out <= 16'h0644;    16'd35461: out <= 16'h067F;    16'd35462: out <= 16'h0195;    16'd35463: out <= 16'h02A6;
    16'd35464: out <= 16'h01E3;    16'd35465: out <= 16'h0538;    16'd35466: out <= 16'h07B2;    16'd35467: out <= 16'h04CA;
    16'd35468: out <= 16'h0ACD;    16'd35469: out <= 16'h0321;    16'd35470: out <= 16'h0447;    16'd35471: out <= 16'h0072;
    16'd35472: out <= 16'h026E;    16'd35473: out <= 16'hFF0B;    16'd35474: out <= 16'h067A;    16'd35475: out <= 16'hFE27;
    16'd35476: out <= 16'h0423;    16'd35477: out <= 16'h07A8;    16'd35478: out <= 16'h04E4;    16'd35479: out <= 16'h003A;
    16'd35480: out <= 16'h057E;    16'd35481: out <= 16'h0592;    16'd35482: out <= 16'h049D;    16'd35483: out <= 16'h0428;
    16'd35484: out <= 16'h0034;    16'd35485: out <= 16'hFBF9;    16'd35486: out <= 16'h030C;    16'd35487: out <= 16'h011A;
    16'd35488: out <= 16'h0A38;    16'd35489: out <= 16'hFBD6;    16'd35490: out <= 16'h0632;    16'd35491: out <= 16'h0C75;
    16'd35492: out <= 16'h092A;    16'd35493: out <= 16'h06AB;    16'd35494: out <= 16'hFC4C;    16'd35495: out <= 16'h03D6;
    16'd35496: out <= 16'hFF41;    16'd35497: out <= 16'h019E;    16'd35498: out <= 16'hFC6C;    16'd35499: out <= 16'h02CF;
    16'd35500: out <= 16'hFEF4;    16'd35501: out <= 16'h0A7E;    16'd35502: out <= 16'hFFFC;    16'd35503: out <= 16'h027E;
    16'd35504: out <= 16'h04B4;    16'd35505: out <= 16'h0530;    16'd35506: out <= 16'h085D;    16'd35507: out <= 16'h0B3F;
    16'd35508: out <= 16'h08D8;    16'd35509: out <= 16'h0623;    16'd35510: out <= 16'hF805;    16'd35511: out <= 16'hFE13;
    16'd35512: out <= 16'h0912;    16'd35513: out <= 16'h072E;    16'd35514: out <= 16'h064F;    16'd35515: out <= 16'h0508;
    16'd35516: out <= 16'h0A04;    16'd35517: out <= 16'h066D;    16'd35518: out <= 16'h09E7;    16'd35519: out <= 16'h0466;
    16'd35520: out <= 16'h0000;    16'd35521: out <= 16'h0652;    16'd35522: out <= 16'h0385;    16'd35523: out <= 16'h023F;
    16'd35524: out <= 16'hFF44;    16'd35525: out <= 16'h03D8;    16'd35526: out <= 16'h0278;    16'd35527: out <= 16'h00AC;
    16'd35528: out <= 16'h017F;    16'd35529: out <= 16'h01BA;    16'd35530: out <= 16'h07B9;    16'd35531: out <= 16'h057B;
    16'd35532: out <= 16'h034E;    16'd35533: out <= 16'h0499;    16'd35534: out <= 16'h0CEE;    16'd35535: out <= 16'hFD2E;
    16'd35536: out <= 16'hFFD4;    16'd35537: out <= 16'hFF43;    16'd35538: out <= 16'h0404;    16'd35539: out <= 16'h0A9B;
    16'd35540: out <= 16'h00F5;    16'd35541: out <= 16'h0678;    16'd35542: out <= 16'h0319;    16'd35543: out <= 16'h019A;
    16'd35544: out <= 16'hFDDF;    16'd35545: out <= 16'h0345;    16'd35546: out <= 16'h0417;    16'd35547: out <= 16'h0351;
    16'd35548: out <= 16'h035B;    16'd35549: out <= 16'h0573;    16'd35550: out <= 16'hFF97;    16'd35551: out <= 16'hFDCC;
    16'd35552: out <= 16'h049C;    16'd35553: out <= 16'h060D;    16'd35554: out <= 16'h08E5;    16'd35555: out <= 16'hFF4A;
    16'd35556: out <= 16'hFD5F;    16'd35557: out <= 16'h09D2;    16'd35558: out <= 16'h03CF;    16'd35559: out <= 16'h0559;
    16'd35560: out <= 16'h0001;    16'd35561: out <= 16'hFDE9;    16'd35562: out <= 16'h0318;    16'd35563: out <= 16'h0081;
    16'd35564: out <= 16'h020B;    16'd35565: out <= 16'hFF76;    16'd35566: out <= 16'hFC5A;    16'd35567: out <= 16'h02D0;
    16'd35568: out <= 16'h008F;    16'd35569: out <= 16'hFEE2;    16'd35570: out <= 16'h0474;    16'd35571: out <= 16'hFAFE;
    16'd35572: out <= 16'hFEDC;    16'd35573: out <= 16'hFECB;    16'd35574: out <= 16'h0177;    16'd35575: out <= 16'hFA74;
    16'd35576: out <= 16'h009B;    16'd35577: out <= 16'hFEB3;    16'd35578: out <= 16'hFB43;    16'd35579: out <= 16'hFD37;
    16'd35580: out <= 16'hFDA0;    16'd35581: out <= 16'h00F8;    16'd35582: out <= 16'hFAD2;    16'd35583: out <= 16'hFBFA;
    16'd35584: out <= 16'hFF7A;    16'd35585: out <= 16'h0941;    16'd35586: out <= 16'h0A87;    16'd35587: out <= 16'hFCD3;
    16'd35588: out <= 16'h0487;    16'd35589: out <= 16'hF795;    16'd35590: out <= 16'h0371;    16'd35591: out <= 16'hFFB7;
    16'd35592: out <= 16'h0264;    16'd35593: out <= 16'hFE08;    16'd35594: out <= 16'h00DC;    16'd35595: out <= 16'hFD5F;
    16'd35596: out <= 16'hFFE6;    16'd35597: out <= 16'h02E1;    16'd35598: out <= 16'h00C9;    16'd35599: out <= 16'hFD77;
    16'd35600: out <= 16'hFCFD;    16'd35601: out <= 16'h02C6;    16'd35602: out <= 16'hFA25;    16'd35603: out <= 16'h036F;
    16'd35604: out <= 16'hFE21;    16'd35605: out <= 16'hFEA8;    16'd35606: out <= 16'hFDFC;    16'd35607: out <= 16'h00C3;
    16'd35608: out <= 16'h0848;    16'd35609: out <= 16'h058A;    16'd35610: out <= 16'h04AB;    16'd35611: out <= 16'h07D8;
    16'd35612: out <= 16'h08AD;    16'd35613: out <= 16'hFFE4;    16'd35614: out <= 16'h0510;    16'd35615: out <= 16'h0E5C;
    16'd35616: out <= 16'h0080;    16'd35617: out <= 16'h080D;    16'd35618: out <= 16'hFE56;    16'd35619: out <= 16'h0344;
    16'd35620: out <= 16'h07C4;    16'd35621: out <= 16'h07EF;    16'd35622: out <= 16'h02D4;    16'd35623: out <= 16'h0490;
    16'd35624: out <= 16'h0622;    16'd35625: out <= 16'h0B87;    16'd35626: out <= 16'h0253;    16'd35627: out <= 16'h0EAE;
    16'd35628: out <= 16'h04FA;    16'd35629: out <= 16'h09D5;    16'd35630: out <= 16'h00CB;    16'd35631: out <= 16'h044E;
    16'd35632: out <= 16'h018A;    16'd35633: out <= 16'hFE66;    16'd35634: out <= 16'h03DE;    16'd35635: out <= 16'h02CE;
    16'd35636: out <= 16'h04D8;    16'd35637: out <= 16'hFEDC;    16'd35638: out <= 16'h05C0;    16'd35639: out <= 16'hFAA1;
    16'd35640: out <= 16'hFDA6;    16'd35641: out <= 16'h0703;    16'd35642: out <= 16'h04BD;    16'd35643: out <= 16'h084A;
    16'd35644: out <= 16'h095B;    16'd35645: out <= 16'h025F;    16'd35646: out <= 16'h05D5;    16'd35647: out <= 16'hFB89;
    16'd35648: out <= 16'h0386;    16'd35649: out <= 16'h09A7;    16'd35650: out <= 16'h0A3F;    16'd35651: out <= 16'h032C;
    16'd35652: out <= 16'h0448;    16'd35653: out <= 16'h01A2;    16'd35654: out <= 16'h06BE;    16'd35655: out <= 16'h05BE;
    16'd35656: out <= 16'h0E57;    16'd35657: out <= 16'h038D;    16'd35658: out <= 16'h0773;    16'd35659: out <= 16'h05D8;
    16'd35660: out <= 16'h093C;    16'd35661: out <= 16'h004F;    16'd35662: out <= 16'h03C1;    16'd35663: out <= 16'hFE4D;
    16'd35664: out <= 16'hFFD5;    16'd35665: out <= 16'h03CA;    16'd35666: out <= 16'h026B;    16'd35667: out <= 16'h037A;
    16'd35668: out <= 16'h051C;    16'd35669: out <= 16'h08F3;    16'd35670: out <= 16'h0072;    16'd35671: out <= 16'h0B25;
    16'd35672: out <= 16'h073C;    16'd35673: out <= 16'h023E;    16'd35674: out <= 16'h0316;    16'd35675: out <= 16'h01F2;
    16'd35676: out <= 16'h040B;    16'd35677: out <= 16'h08A4;    16'd35678: out <= 16'h0D70;    16'd35679: out <= 16'hFCAD;
    16'd35680: out <= 16'h0193;    16'd35681: out <= 16'h0490;    16'd35682: out <= 16'h0801;    16'd35683: out <= 16'h0390;
    16'd35684: out <= 16'h042B;    16'd35685: out <= 16'h007B;    16'd35686: out <= 16'h006E;    16'd35687: out <= 16'h0A51;
    16'd35688: out <= 16'h0D71;    16'd35689: out <= 16'h0337;    16'd35690: out <= 16'h05F8;    16'd35691: out <= 16'h0899;
    16'd35692: out <= 16'h0559;    16'd35693: out <= 16'h0487;    16'd35694: out <= 16'h012B;    16'd35695: out <= 16'h03D5;
    16'd35696: out <= 16'h013A;    16'd35697: out <= 16'h03BA;    16'd35698: out <= 16'h0258;    16'd35699: out <= 16'h017A;
    16'd35700: out <= 16'h05A1;    16'd35701: out <= 16'h0777;    16'd35702: out <= 16'h095C;    16'd35703: out <= 16'h0047;
    16'd35704: out <= 16'h01BB;    16'd35705: out <= 16'hFBA2;    16'd35706: out <= 16'h08DA;    16'd35707: out <= 16'hFF26;
    16'd35708: out <= 16'hFECA;    16'd35709: out <= 16'h05AD;    16'd35710: out <= 16'h07FF;    16'd35711: out <= 16'hFE25;
    16'd35712: out <= 16'h024F;    16'd35713: out <= 16'h024E;    16'd35714: out <= 16'h0CBF;    16'd35715: out <= 16'h00A8;
    16'd35716: out <= 16'h0508;    16'd35717: out <= 16'h017C;    16'd35718: out <= 16'h01AC;    16'd35719: out <= 16'h02FB;
    16'd35720: out <= 16'h0E36;    16'd35721: out <= 16'hFE67;    16'd35722: out <= 16'h0BA2;    16'd35723: out <= 16'h0543;
    16'd35724: out <= 16'h0BF6;    16'd35725: out <= 16'h0190;    16'd35726: out <= 16'hFD44;    16'd35727: out <= 16'h0263;
    16'd35728: out <= 16'h00BA;    16'd35729: out <= 16'h0765;    16'd35730: out <= 16'h006D;    16'd35731: out <= 16'h0687;
    16'd35732: out <= 16'h0253;    16'd35733: out <= 16'h0333;    16'd35734: out <= 16'h09F7;    16'd35735: out <= 16'h0371;
    16'd35736: out <= 16'h0166;    16'd35737: out <= 16'h0497;    16'd35738: out <= 16'h07B1;    16'd35739: out <= 16'hFFC9;
    16'd35740: out <= 16'h00C9;    16'd35741: out <= 16'hFF8B;    16'd35742: out <= 16'h0534;    16'd35743: out <= 16'h09A3;
    16'd35744: out <= 16'hFFD8;    16'd35745: out <= 16'h01DB;    16'd35746: out <= 16'h0C7E;    16'd35747: out <= 16'hFEDC;
    16'd35748: out <= 16'h0574;    16'd35749: out <= 16'h0A7E;    16'd35750: out <= 16'h0718;    16'd35751: out <= 16'h053A;
    16'd35752: out <= 16'h0CE3;    16'd35753: out <= 16'h0266;    16'd35754: out <= 16'h0488;    16'd35755: out <= 16'h0690;
    16'd35756: out <= 16'h06DE;    16'd35757: out <= 16'h03CA;    16'd35758: out <= 16'hFD27;    16'd35759: out <= 16'h040B;
    16'd35760: out <= 16'h01DA;    16'd35761: out <= 16'h0537;    16'd35762: out <= 16'h01AC;    16'd35763: out <= 16'h029A;
    16'd35764: out <= 16'h01B4;    16'd35765: out <= 16'h062E;    16'd35766: out <= 16'h06A8;    16'd35767: out <= 16'h02CD;
    16'd35768: out <= 16'h00CA;    16'd35769: out <= 16'h04F6;    16'd35770: out <= 16'hFF12;    16'd35771: out <= 16'hFF6F;
    16'd35772: out <= 16'h0769;    16'd35773: out <= 16'h0846;    16'd35774: out <= 16'h0357;    16'd35775: out <= 16'h050B;
    16'd35776: out <= 16'h00E2;    16'd35777: out <= 16'hFF36;    16'd35778: out <= 16'h03D3;    16'd35779: out <= 16'h0971;
    16'd35780: out <= 16'h039E;    16'd35781: out <= 16'h0807;    16'd35782: out <= 16'h0877;    16'd35783: out <= 16'h0732;
    16'd35784: out <= 16'h027F;    16'd35785: out <= 16'h01EB;    16'd35786: out <= 16'hF94A;    16'd35787: out <= 16'h0489;
    16'd35788: out <= 16'h06C1;    16'd35789: out <= 16'h0239;    16'd35790: out <= 16'h022F;    16'd35791: out <= 16'h09C9;
    16'd35792: out <= 16'h09E6;    16'd35793: out <= 16'h06D6;    16'd35794: out <= 16'h08A0;    16'd35795: out <= 16'h0265;
    16'd35796: out <= 16'h0649;    16'd35797: out <= 16'h02F5;    16'd35798: out <= 16'h02A1;    16'd35799: out <= 16'h0333;
    16'd35800: out <= 16'h0154;    16'd35801: out <= 16'hFD3B;    16'd35802: out <= 16'h0079;    16'd35803: out <= 16'h015D;
    16'd35804: out <= 16'h0544;    16'd35805: out <= 16'h08E9;    16'd35806: out <= 16'h07DE;    16'd35807: out <= 16'h044C;
    16'd35808: out <= 16'h0676;    16'd35809: out <= 16'h014E;    16'd35810: out <= 16'h016B;    16'd35811: out <= 16'h012A;
    16'd35812: out <= 16'h0A87;    16'd35813: out <= 16'h038F;    16'd35814: out <= 16'hFDF4;    16'd35815: out <= 16'h05F5;
    16'd35816: out <= 16'h01B2;    16'd35817: out <= 16'h007D;    16'd35818: out <= 16'h0221;    16'd35819: out <= 16'h031C;
    16'd35820: out <= 16'hFDB4;    16'd35821: out <= 16'h082A;    16'd35822: out <= 16'h03FF;    16'd35823: out <= 16'h033B;
    16'd35824: out <= 16'hFD4D;    16'd35825: out <= 16'h01CD;    16'd35826: out <= 16'h05AE;    16'd35827: out <= 16'hFE16;
    16'd35828: out <= 16'hFDA6;    16'd35829: out <= 16'hFFA1;    16'd35830: out <= 16'hFFD2;    16'd35831: out <= 16'hFDDF;
    16'd35832: out <= 16'h0734;    16'd35833: out <= 16'hFA2B;    16'd35834: out <= 16'h04AB;    16'd35835: out <= 16'h00F2;
    16'd35836: out <= 16'hFF44;    16'd35837: out <= 16'hFB86;    16'd35838: out <= 16'h0756;    16'd35839: out <= 16'hF812;
    16'd35840: out <= 16'hF72B;    16'd35841: out <= 16'hFB69;    16'd35842: out <= 16'h053B;    16'd35843: out <= 16'h009E;
    16'd35844: out <= 16'hF8A5;    16'd35845: out <= 16'h02B2;    16'd35846: out <= 16'hF753;    16'd35847: out <= 16'h0398;
    16'd35848: out <= 16'hFC77;    16'd35849: out <= 16'h0180;    16'd35850: out <= 16'hFF8D;    16'd35851: out <= 16'hFFE3;
    16'd35852: out <= 16'hFD77;    16'd35853: out <= 16'hFF99;    16'd35854: out <= 16'h00E4;    16'd35855: out <= 16'hF8EB;
    16'd35856: out <= 16'hFAC0;    16'd35857: out <= 16'h0475;    16'd35858: out <= 16'h07F1;    16'd35859: out <= 16'h022E;
    16'd35860: out <= 16'h00CD;    16'd35861: out <= 16'h0405;    16'd35862: out <= 16'h034C;    16'd35863: out <= 16'hFE12;
    16'd35864: out <= 16'h049A;    16'd35865: out <= 16'h0884;    16'd35866: out <= 16'h0DCC;    16'd35867: out <= 16'hF91C;
    16'd35868: out <= 16'h0168;    16'd35869: out <= 16'h04BD;    16'd35870: out <= 16'hFDA8;    16'd35871: out <= 16'h0488;
    16'd35872: out <= 16'hFC7E;    16'd35873: out <= 16'h0468;    16'd35874: out <= 16'hFBF0;    16'd35875: out <= 16'hFEB8;
    16'd35876: out <= 16'h0AE7;    16'd35877: out <= 16'h0012;    16'd35878: out <= 16'h00E7;    16'd35879: out <= 16'h047F;
    16'd35880: out <= 16'h0247;    16'd35881: out <= 16'h0306;    16'd35882: out <= 16'hFF2E;    16'd35883: out <= 16'hFFB4;
    16'd35884: out <= 16'h0478;    16'd35885: out <= 16'hFDB7;    16'd35886: out <= 16'h0327;    16'd35887: out <= 16'h0536;
    16'd35888: out <= 16'h04B8;    16'd35889: out <= 16'h0386;    16'd35890: out <= 16'hFD72;    16'd35891: out <= 16'h01D6;
    16'd35892: out <= 16'h0732;    16'd35893: out <= 16'h05B4;    16'd35894: out <= 16'h08D7;    16'd35895: out <= 16'h005D;
    16'd35896: out <= 16'hFFD2;    16'd35897: out <= 16'h0234;    16'd35898: out <= 16'h02DB;    16'd35899: out <= 16'h045E;
    16'd35900: out <= 16'h0263;    16'd35901: out <= 16'hFFEB;    16'd35902: out <= 16'h0828;    16'd35903: out <= 16'h01AC;
    16'd35904: out <= 16'h045D;    16'd35905: out <= 16'h0959;    16'd35906: out <= 16'h0152;    16'd35907: out <= 16'h0419;
    16'd35908: out <= 16'h00B1;    16'd35909: out <= 16'hFC3B;    16'd35910: out <= 16'hFFE2;    16'd35911: out <= 16'h0501;
    16'd35912: out <= 16'h052B;    16'd35913: out <= 16'hFF60;    16'd35914: out <= 16'h0529;    16'd35915: out <= 16'h029F;
    16'd35916: out <= 16'h0059;    16'd35917: out <= 16'h05E8;    16'd35918: out <= 16'h02BB;    16'd35919: out <= 16'h0875;
    16'd35920: out <= 16'h0580;    16'd35921: out <= 16'h0301;    16'd35922: out <= 16'h01CF;    16'd35923: out <= 16'h074B;
    16'd35924: out <= 16'h0214;    16'd35925: out <= 16'h01DC;    16'd35926: out <= 16'hFD85;    16'd35927: out <= 16'hFCEB;
    16'd35928: out <= 16'hFFEC;    16'd35929: out <= 16'h021A;    16'd35930: out <= 16'h01D1;    16'd35931: out <= 16'h00BE;
    16'd35932: out <= 16'h00E0;    16'd35933: out <= 16'h0701;    16'd35934: out <= 16'h006A;    16'd35935: out <= 16'hFD1E;
    16'd35936: out <= 16'h057C;    16'd35937: out <= 16'h07BD;    16'd35938: out <= 16'h008F;    16'd35939: out <= 16'h07E5;
    16'd35940: out <= 16'h0186;    16'd35941: out <= 16'h0AE7;    16'd35942: out <= 16'h02E9;    16'd35943: out <= 16'hFD88;
    16'd35944: out <= 16'hFFCD;    16'd35945: out <= 16'h0155;    16'd35946: out <= 16'h0368;    16'd35947: out <= 16'hFD3D;
    16'd35948: out <= 16'h064B;    16'd35949: out <= 16'hFF55;    16'd35950: out <= 16'h06BB;    16'd35951: out <= 16'h02E7;
    16'd35952: out <= 16'h061A;    16'd35953: out <= 16'h0477;    16'd35954: out <= 16'h0821;    16'd35955: out <= 16'h04E8;
    16'd35956: out <= 16'h04B3;    16'd35957: out <= 16'h0704;    16'd35958: out <= 16'h042F;    16'd35959: out <= 16'h080B;
    16'd35960: out <= 16'h02CC;    16'd35961: out <= 16'h0B87;    16'd35962: out <= 16'h00B9;    16'd35963: out <= 16'h0B89;
    16'd35964: out <= 16'h0056;    16'd35965: out <= 16'h037D;    16'd35966: out <= 16'h01B1;    16'd35967: out <= 16'h01E6;
    16'd35968: out <= 16'h0A99;    16'd35969: out <= 16'h02A8;    16'd35970: out <= 16'hFF75;    16'd35971: out <= 16'h01DD;
    16'd35972: out <= 16'h0287;    16'd35973: out <= 16'h0208;    16'd35974: out <= 16'h0411;    16'd35975: out <= 16'hF833;
    16'd35976: out <= 16'hFDC3;    16'd35977: out <= 16'h0239;    16'd35978: out <= 16'h02B8;    16'd35979: out <= 16'h05BB;
    16'd35980: out <= 16'h02DB;    16'd35981: out <= 16'h04E8;    16'd35982: out <= 16'h0B01;    16'd35983: out <= 16'h04A2;
    16'd35984: out <= 16'hFF40;    16'd35985: out <= 16'hFFA4;    16'd35986: out <= 16'h089A;    16'd35987: out <= 16'h0BFD;
    16'd35988: out <= 16'h0472;    16'd35989: out <= 16'h026D;    16'd35990: out <= 16'h0109;    16'd35991: out <= 16'h0225;
    16'd35992: out <= 16'h0503;    16'd35993: out <= 16'h0708;    16'd35994: out <= 16'h036F;    16'd35995: out <= 16'h035A;
    16'd35996: out <= 16'hFE67;    16'd35997: out <= 16'h04FD;    16'd35998: out <= 16'h05BC;    16'd35999: out <= 16'h02C1;
    16'd36000: out <= 16'h076B;    16'd36001: out <= 16'hFCEC;    16'd36002: out <= 16'hFC5B;    16'd36003: out <= 16'h0009;
    16'd36004: out <= 16'h00B2;    16'd36005: out <= 16'h0314;    16'd36006: out <= 16'h0748;    16'd36007: out <= 16'h074E;
    16'd36008: out <= 16'h0814;    16'd36009: out <= 16'h04FB;    16'd36010: out <= 16'h06CA;    16'd36011: out <= 16'h0485;
    16'd36012: out <= 16'h02CF;    16'd36013: out <= 16'h012D;    16'd36014: out <= 16'h0802;    16'd36015: out <= 16'h04DE;
    16'd36016: out <= 16'h046D;    16'd36017: out <= 16'h028C;    16'd36018: out <= 16'h0331;    16'd36019: out <= 16'h04DD;
    16'd36020: out <= 16'h06F4;    16'd36021: out <= 16'hFE12;    16'd36022: out <= 16'h005D;    16'd36023: out <= 16'h05F5;
    16'd36024: out <= 16'h0A19;    16'd36025: out <= 16'h0A10;    16'd36026: out <= 16'h02C4;    16'd36027: out <= 16'hF768;
    16'd36028: out <= 16'h003A;    16'd36029: out <= 16'h064D;    16'd36030: out <= 16'h007C;    16'd36031: out <= 16'h0648;
    16'd36032: out <= 16'h039D;    16'd36033: out <= 16'h051A;    16'd36034: out <= 16'h056B;    16'd36035: out <= 16'h02B2;
    16'd36036: out <= 16'h0516;    16'd36037: out <= 16'h00C7;    16'd36038: out <= 16'hFF52;    16'd36039: out <= 16'h060C;
    16'd36040: out <= 16'h0A8E;    16'd36041: out <= 16'h0700;    16'd36042: out <= 16'h03DD;    16'd36043: out <= 16'h0469;
    16'd36044: out <= 16'h027F;    16'd36045: out <= 16'hFDF2;    16'd36046: out <= 16'h025D;    16'd36047: out <= 16'h046E;
    16'd36048: out <= 16'h02D0;    16'd36049: out <= 16'h04CD;    16'd36050: out <= 16'h08CA;    16'd36051: out <= 16'h07E1;
    16'd36052: out <= 16'h03B6;    16'd36053: out <= 16'h0004;    16'd36054: out <= 16'h0C16;    16'd36055: out <= 16'h080F;
    16'd36056: out <= 16'hFDC3;    16'd36057: out <= 16'hFEC9;    16'd36058: out <= 16'h039D;    16'd36059: out <= 16'h0068;
    16'd36060: out <= 16'hFFE7;    16'd36061: out <= 16'h0C73;    16'd36062: out <= 16'h00B4;    16'd36063: out <= 16'h0412;
    16'd36064: out <= 16'h0420;    16'd36065: out <= 16'h04D0;    16'd36066: out <= 16'hFF19;    16'd36067: out <= 16'h072A;
    16'd36068: out <= 16'h03EB;    16'd36069: out <= 16'h04B4;    16'd36070: out <= 16'h083F;    16'd36071: out <= 16'h0437;
    16'd36072: out <= 16'hFF61;    16'd36073: out <= 16'hFE0C;    16'd36074: out <= 16'hFD23;    16'd36075: out <= 16'hFDDB;
    16'd36076: out <= 16'hFB00;    16'd36077: out <= 16'h0065;    16'd36078: out <= 16'h008A;    16'd36079: out <= 16'hFE63;
    16'd36080: out <= 16'h0134;    16'd36081: out <= 16'hFB34;    16'd36082: out <= 16'h02F3;    16'd36083: out <= 16'hFBE9;
    16'd36084: out <= 16'h037F;    16'd36085: out <= 16'h0532;    16'd36086: out <= 16'hFE47;    16'd36087: out <= 16'h0330;
    16'd36088: out <= 16'hFCB7;    16'd36089: out <= 16'h0100;    16'd36090: out <= 16'hFDD0;    16'd36091: out <= 16'hFDCB;
    16'd36092: out <= 16'hFCEF;    16'd36093: out <= 16'hFA89;    16'd36094: out <= 16'hFC9F;    16'd36095: out <= 16'h02D7;
    16'd36096: out <= 16'hFA93;    16'd36097: out <= 16'h0261;    16'd36098: out <= 16'hFFBD;    16'd36099: out <= 16'hFE57;
    16'd36100: out <= 16'h02FD;    16'd36101: out <= 16'h031E;    16'd36102: out <= 16'h0488;    16'd36103: out <= 16'h0560;
    16'd36104: out <= 16'h01B8;    16'd36105: out <= 16'hFED5;    16'd36106: out <= 16'hFE38;    16'd36107: out <= 16'h0668;
    16'd36108: out <= 16'h01B7;    16'd36109: out <= 16'hFBB4;    16'd36110: out <= 16'hFDAE;    16'd36111: out <= 16'hFEEB;
    16'd36112: out <= 16'h02F9;    16'd36113: out <= 16'h02E7;    16'd36114: out <= 16'hFFFC;    16'd36115: out <= 16'h0048;
    16'd36116: out <= 16'h06F6;    16'd36117: out <= 16'hFA13;    16'd36118: out <= 16'hF8CF;    16'd36119: out <= 16'h035C;
    16'd36120: out <= 16'h05A0;    16'd36121: out <= 16'h000E;    16'd36122: out <= 16'hFECC;    16'd36123: out <= 16'hFFA2;
    16'd36124: out <= 16'h0227;    16'd36125: out <= 16'hFE87;    16'd36126: out <= 16'h03EC;    16'd36127: out <= 16'h00B9;
    16'd36128: out <= 16'h02AF;    16'd36129: out <= 16'hFDBB;    16'd36130: out <= 16'h0B04;    16'd36131: out <= 16'h0514;
    16'd36132: out <= 16'h0600;    16'd36133: out <= 16'h0416;    16'd36134: out <= 16'h00B5;    16'd36135: out <= 16'h05B8;
    16'd36136: out <= 16'h0C07;    16'd36137: out <= 16'h02AB;    16'd36138: out <= 16'hFA65;    16'd36139: out <= 16'h0C3B;
    16'd36140: out <= 16'h05D0;    16'd36141: out <= 16'h05EC;    16'd36142: out <= 16'h0598;    16'd36143: out <= 16'h0143;
    16'd36144: out <= 16'hFBBF;    16'd36145: out <= 16'h0C64;    16'd36146: out <= 16'h0B01;    16'd36147: out <= 16'h01B8;
    16'd36148: out <= 16'h0496;    16'd36149: out <= 16'h06CD;    16'd36150: out <= 16'hFDB5;    16'd36151: out <= 16'h0216;
    16'd36152: out <= 16'h0628;    16'd36153: out <= 16'hFE64;    16'd36154: out <= 16'h084F;    16'd36155: out <= 16'h0312;
    16'd36156: out <= 16'h050E;    16'd36157: out <= 16'h0774;    16'd36158: out <= 16'h03DE;    16'd36159: out <= 16'h0772;
    16'd36160: out <= 16'h072D;    16'd36161: out <= 16'hFDC0;    16'd36162: out <= 16'h00FF;    16'd36163: out <= 16'h0282;
    16'd36164: out <= 16'h07B6;    16'd36165: out <= 16'h0353;    16'd36166: out <= 16'h0314;    16'd36167: out <= 16'hFF34;
    16'd36168: out <= 16'h0E97;    16'd36169: out <= 16'h088D;    16'd36170: out <= 16'h0254;    16'd36171: out <= 16'hFEFC;
    16'd36172: out <= 16'h05C3;    16'd36173: out <= 16'h0304;    16'd36174: out <= 16'h0F64;    16'd36175: out <= 16'h01F2;
    16'd36176: out <= 16'h0383;    16'd36177: out <= 16'h04D5;    16'd36178: out <= 16'h00FD;    16'd36179: out <= 16'hFF18;
    16'd36180: out <= 16'h0218;    16'd36181: out <= 16'h0452;    16'd36182: out <= 16'h0B2E;    16'd36183: out <= 16'h0BD3;
    16'd36184: out <= 16'h016D;    16'd36185: out <= 16'h042E;    16'd36186: out <= 16'h0694;    16'd36187: out <= 16'h0457;
    16'd36188: out <= 16'h0314;    16'd36189: out <= 16'h05BA;    16'd36190: out <= 16'h01C6;    16'd36191: out <= 16'h0A2A;
    16'd36192: out <= 16'h020D;    16'd36193: out <= 16'h046B;    16'd36194: out <= 16'h03F2;    16'd36195: out <= 16'h031B;
    16'd36196: out <= 16'h0459;    16'd36197: out <= 16'hFDB7;    16'd36198: out <= 16'hFF47;    16'd36199: out <= 16'hFDAC;
    16'd36200: out <= 16'h00CB;    16'd36201: out <= 16'h0519;    16'd36202: out <= 16'h0568;    16'd36203: out <= 16'h05C3;
    16'd36204: out <= 16'h07C0;    16'd36205: out <= 16'h0231;    16'd36206: out <= 16'h08D5;    16'd36207: out <= 16'h0575;
    16'd36208: out <= 16'hFF08;    16'd36209: out <= 16'h0967;    16'd36210: out <= 16'hFF89;    16'd36211: out <= 16'hFD54;
    16'd36212: out <= 16'h02FB;    16'd36213: out <= 16'h065D;    16'd36214: out <= 16'h07CD;    16'd36215: out <= 16'h0136;
    16'd36216: out <= 16'h0229;    16'd36217: out <= 16'h030B;    16'd36218: out <= 16'h0793;    16'd36219: out <= 16'h07CF;
    16'd36220: out <= 16'h037B;    16'd36221: out <= 16'hFEDC;    16'd36222: out <= 16'h0AD4;    16'd36223: out <= 16'h062E;
    16'd36224: out <= 16'h0800;    16'd36225: out <= 16'h034C;    16'd36226: out <= 16'h043F;    16'd36227: out <= 16'hFE1D;
    16'd36228: out <= 16'hFF7B;    16'd36229: out <= 16'hFF74;    16'd36230: out <= 16'h06E1;    16'd36231: out <= 16'hFD5E;
    16'd36232: out <= 16'hFFDA;    16'd36233: out <= 16'h08AC;    16'd36234: out <= 16'hFFE8;    16'd36235: out <= 16'h0466;
    16'd36236: out <= 16'h0302;    16'd36237: out <= 16'hFFFF;    16'd36238: out <= 16'h05B1;    16'd36239: out <= 16'hFEE6;
    16'd36240: out <= 16'h016E;    16'd36241: out <= 16'hFD69;    16'd36242: out <= 16'h01AA;    16'd36243: out <= 16'h07CD;
    16'd36244: out <= 16'h077A;    16'd36245: out <= 16'h0170;    16'd36246: out <= 16'h0810;    16'd36247: out <= 16'h0575;
    16'd36248: out <= 16'h083B;    16'd36249: out <= 16'h0894;    16'd36250: out <= 16'h09B0;    16'd36251: out <= 16'h03DE;
    16'd36252: out <= 16'h05C6;    16'd36253: out <= 16'hFCDB;    16'd36254: out <= 16'h04AF;    16'd36255: out <= 16'h028F;
    16'd36256: out <= 16'h01DC;    16'd36257: out <= 16'h0898;    16'd36258: out <= 16'h043E;    16'd36259: out <= 16'h0572;
    16'd36260: out <= 16'h0703;    16'd36261: out <= 16'h085C;    16'd36262: out <= 16'h0650;    16'd36263: out <= 16'h016E;
    16'd36264: out <= 16'h08B1;    16'd36265: out <= 16'h0BB0;    16'd36266: out <= 16'h0621;    16'd36267: out <= 16'h0971;
    16'd36268: out <= 16'hFB3C;    16'd36269: out <= 16'h0AD2;    16'd36270: out <= 16'h0B75;    16'd36271: out <= 16'h0739;
    16'd36272: out <= 16'h02D5;    16'd36273: out <= 16'h039E;    16'd36274: out <= 16'h086C;    16'd36275: out <= 16'h0129;
    16'd36276: out <= 16'h0712;    16'd36277: out <= 16'h056F;    16'd36278: out <= 16'h06A8;    16'd36279: out <= 16'h075A;
    16'd36280: out <= 16'h0028;    16'd36281: out <= 16'hFE6B;    16'd36282: out <= 16'hFA46;    16'd36283: out <= 16'h0371;
    16'd36284: out <= 16'h0C1E;    16'd36285: out <= 16'h0289;    16'd36286: out <= 16'hFE10;    16'd36287: out <= 16'hFE4E;
    16'd36288: out <= 16'h0529;    16'd36289: out <= 16'h04EE;    16'd36290: out <= 16'h0C93;    16'd36291: out <= 16'h007E;
    16'd36292: out <= 16'h0570;    16'd36293: out <= 16'h062D;    16'd36294: out <= 16'h0035;    16'd36295: out <= 16'h0617;
    16'd36296: out <= 16'h0563;    16'd36297: out <= 16'h05FF;    16'd36298: out <= 16'h0568;    16'd36299: out <= 16'hFFF9;
    16'd36300: out <= 16'hFF91;    16'd36301: out <= 16'h0327;    16'd36302: out <= 16'h0950;    16'd36303: out <= 16'hFEFE;
    16'd36304: out <= 16'hFF3B;    16'd36305: out <= 16'h0437;    16'd36306: out <= 16'h0E6B;    16'd36307: out <= 16'h063A;
    16'd36308: out <= 16'hFC99;    16'd36309: out <= 16'hFE81;    16'd36310: out <= 16'hF9F0;    16'd36311: out <= 16'h07CC;
    16'd36312: out <= 16'hF9CB;    16'd36313: out <= 16'hFB24;    16'd36314: out <= 16'hFC19;    16'd36315: out <= 16'h09A7;
    16'd36316: out <= 16'h09D1;    16'd36317: out <= 16'h06EC;    16'd36318: out <= 16'h05C5;    16'd36319: out <= 16'hFE4E;
    16'd36320: out <= 16'h0886;    16'd36321: out <= 16'h0963;    16'd36322: out <= 16'hFEAD;    16'd36323: out <= 16'h0AEA;
    16'd36324: out <= 16'hFB66;    16'd36325: out <= 16'h0210;    16'd36326: out <= 16'h1019;    16'd36327: out <= 16'h087A;
    16'd36328: out <= 16'h04D6;    16'd36329: out <= 16'h07F9;    16'd36330: out <= 16'hFDEC;    16'd36331: out <= 16'hFCAA;
    16'd36332: out <= 16'h0098;    16'd36333: out <= 16'h0338;    16'd36334: out <= 16'h0465;    16'd36335: out <= 16'hF5E8;
    16'd36336: out <= 16'h03A2;    16'd36337: out <= 16'hFC83;    16'd36338: out <= 16'hFC97;    16'd36339: out <= 16'hFD95;
    16'd36340: out <= 16'hFF2F;    16'd36341: out <= 16'hFF41;    16'd36342: out <= 16'h069E;    16'd36343: out <= 16'h015E;
    16'd36344: out <= 16'hFEF6;    16'd36345: out <= 16'hFFB6;    16'd36346: out <= 16'hFC02;    16'd36347: out <= 16'h02FE;
    16'd36348: out <= 16'hFEA4;    16'd36349: out <= 16'h0095;    16'd36350: out <= 16'h00D7;    16'd36351: out <= 16'h082E;
    16'd36352: out <= 16'h021D;    16'd36353: out <= 16'hFEE3;    16'd36354: out <= 16'h0710;    16'd36355: out <= 16'hF897;
    16'd36356: out <= 16'h028C;    16'd36357: out <= 16'h0914;    16'd36358: out <= 16'hFE94;    16'd36359: out <= 16'h0064;
    16'd36360: out <= 16'hFE19;    16'd36361: out <= 16'h0045;    16'd36362: out <= 16'hF6BC;    16'd36363: out <= 16'hFC2F;
    16'd36364: out <= 16'hFB10;    16'd36365: out <= 16'hFB39;    16'd36366: out <= 16'hFDE1;    16'd36367: out <= 16'h00F4;
    16'd36368: out <= 16'hFB68;    16'd36369: out <= 16'h01B8;    16'd36370: out <= 16'h064D;    16'd36371: out <= 16'hFE6A;
    16'd36372: out <= 16'h01C6;    16'd36373: out <= 16'h0012;    16'd36374: out <= 16'hFD42;    16'd36375: out <= 16'h0009;
    16'd36376: out <= 16'hFBEA;    16'd36377: out <= 16'h0576;    16'd36378: out <= 16'h050A;    16'd36379: out <= 16'h096A;
    16'd36380: out <= 16'h0932;    16'd36381: out <= 16'h063C;    16'd36382: out <= 16'h04B3;    16'd36383: out <= 16'h02A2;
    16'd36384: out <= 16'hFFF1;    16'd36385: out <= 16'h050D;    16'd36386: out <= 16'h028D;    16'd36387: out <= 16'h0715;
    16'd36388: out <= 16'h0264;    16'd36389: out <= 16'hFEED;    16'd36390: out <= 16'h0A41;    16'd36391: out <= 16'h0B19;
    16'd36392: out <= 16'h044A;    16'd36393: out <= 16'h090C;    16'd36394: out <= 16'h06C0;    16'd36395: out <= 16'hFEA4;
    16'd36396: out <= 16'hFE47;    16'd36397: out <= 16'h08D2;    16'd36398: out <= 16'hFEB0;    16'd36399: out <= 16'h01B8;
    16'd36400: out <= 16'h0438;    16'd36401: out <= 16'hFE4D;    16'd36402: out <= 16'h0386;    16'd36403: out <= 16'h00D1;
    16'd36404: out <= 16'h0540;    16'd36405: out <= 16'h050C;    16'd36406: out <= 16'hFEC8;    16'd36407: out <= 16'h04FE;
    16'd36408: out <= 16'h0377;    16'd36409: out <= 16'h00DF;    16'd36410: out <= 16'hFFB7;    16'd36411: out <= 16'h07C6;
    16'd36412: out <= 16'h0D21;    16'd36413: out <= 16'hFEAA;    16'd36414: out <= 16'h08EC;    16'd36415: out <= 16'hFFFD;
    16'd36416: out <= 16'h0BAA;    16'd36417: out <= 16'h03E4;    16'd36418: out <= 16'h063D;    16'd36419: out <= 16'hFCA4;
    16'd36420: out <= 16'h04F1;    16'd36421: out <= 16'h00DF;    16'd36422: out <= 16'h00CB;    16'd36423: out <= 16'h001F;
    16'd36424: out <= 16'hFEC9;    16'd36425: out <= 16'h04A6;    16'd36426: out <= 16'h0555;    16'd36427: out <= 16'hFD1E;
    16'd36428: out <= 16'hFDB9;    16'd36429: out <= 16'h09DE;    16'd36430: out <= 16'h0552;    16'd36431: out <= 16'h05DD;
    16'd36432: out <= 16'h0665;    16'd36433: out <= 16'h05AF;    16'd36434: out <= 16'h033F;    16'd36435: out <= 16'h01D9;
    16'd36436: out <= 16'h00AF;    16'd36437: out <= 16'h02D0;    16'd36438: out <= 16'h02B4;    16'd36439: out <= 16'hFF8F;
    16'd36440: out <= 16'h08A1;    16'd36441: out <= 16'h07AB;    16'd36442: out <= 16'hFB33;    16'd36443: out <= 16'hFED7;
    16'd36444: out <= 16'hFC43;    16'd36445: out <= 16'h0606;    16'd36446: out <= 16'h05FF;    16'd36447: out <= 16'h04E2;
    16'd36448: out <= 16'h04C2;    16'd36449: out <= 16'h0205;    16'd36450: out <= 16'h03B9;    16'd36451: out <= 16'h0608;
    16'd36452: out <= 16'h03BC;    16'd36453: out <= 16'hFCAC;    16'd36454: out <= 16'h044E;    16'd36455: out <= 16'hF786;
    16'd36456: out <= 16'hFF83;    16'd36457: out <= 16'hFBC4;    16'd36458: out <= 16'hFE4A;    16'd36459: out <= 16'h03A1;
    16'd36460: out <= 16'h060F;    16'd36461: out <= 16'hFEE2;    16'd36462: out <= 16'h065C;    16'd36463: out <= 16'h0A11;
    16'd36464: out <= 16'h0133;    16'd36465: out <= 16'h02D9;    16'd36466: out <= 16'hFD50;    16'd36467: out <= 16'h0303;
    16'd36468: out <= 16'hFCED;    16'd36469: out <= 16'h00A4;    16'd36470: out <= 16'hFEB6;    16'd36471: out <= 16'hFE8B;
    16'd36472: out <= 16'h0811;    16'd36473: out <= 16'h0624;    16'd36474: out <= 16'h09E4;    16'd36475: out <= 16'hFF82;
    16'd36476: out <= 16'h004D;    16'd36477: out <= 16'h044E;    16'd36478: out <= 16'h0202;    16'd36479: out <= 16'h0080;
    16'd36480: out <= 16'h001F;    16'd36481: out <= 16'h0031;    16'd36482: out <= 16'h0429;    16'd36483: out <= 16'hFAD8;
    16'd36484: out <= 16'h03CE;    16'd36485: out <= 16'hFE78;    16'd36486: out <= 16'hFD96;    16'd36487: out <= 16'h00BF;
    16'd36488: out <= 16'hFC5D;    16'd36489: out <= 16'h00C9;    16'd36490: out <= 16'h0287;    16'd36491: out <= 16'h054F;
    16'd36492: out <= 16'h0198;    16'd36493: out <= 16'h0653;    16'd36494: out <= 16'h0122;    16'd36495: out <= 16'hFF47;
    16'd36496: out <= 16'h02F6;    16'd36497: out <= 16'h021B;    16'd36498: out <= 16'hFF5D;    16'd36499: out <= 16'hFCA7;
    16'd36500: out <= 16'h08C4;    16'd36501: out <= 16'h0000;    16'd36502: out <= 16'h086F;    16'd36503: out <= 16'h0962;
    16'd36504: out <= 16'hFF9A;    16'd36505: out <= 16'h03DC;    16'd36506: out <= 16'h031D;    16'd36507: out <= 16'h0043;
    16'd36508: out <= 16'h0547;    16'd36509: out <= 16'h01E6;    16'd36510: out <= 16'h063F;    16'd36511: out <= 16'h0AA9;
    16'd36512: out <= 16'h0533;    16'd36513: out <= 16'hFBD9;    16'd36514: out <= 16'hFF90;    16'd36515: out <= 16'h02FF;
    16'd36516: out <= 16'h01EA;    16'd36517: out <= 16'hFFF3;    16'd36518: out <= 16'h08C6;    16'd36519: out <= 16'h00DB;
    16'd36520: out <= 16'h0102;    16'd36521: out <= 16'h0466;    16'd36522: out <= 16'h07C1;    16'd36523: out <= 16'hFF85;
    16'd36524: out <= 16'h06D0;    16'd36525: out <= 16'h003F;    16'd36526: out <= 16'hFF00;    16'd36527: out <= 16'h0534;
    16'd36528: out <= 16'h0122;    16'd36529: out <= 16'h083F;    16'd36530: out <= 16'h0922;    16'd36531: out <= 16'h0671;
    16'd36532: out <= 16'h03EA;    16'd36533: out <= 16'h08BE;    16'd36534: out <= 16'h02DB;    16'd36535: out <= 16'h0418;
    16'd36536: out <= 16'h007F;    16'd36537: out <= 16'hFD8F;    16'd36538: out <= 16'h0815;    16'd36539: out <= 16'h062A;
    16'd36540: out <= 16'h00B0;    16'd36541: out <= 16'h0695;    16'd36542: out <= 16'h0527;    16'd36543: out <= 16'h0111;
    16'd36544: out <= 16'hFED9;    16'd36545: out <= 16'h08F7;    16'd36546: out <= 16'hFB44;    16'd36547: out <= 16'hFF7A;
    16'd36548: out <= 16'h0B3E;    16'd36549: out <= 16'h02E9;    16'd36550: out <= 16'h0401;    16'd36551: out <= 16'hFC7E;
    16'd36552: out <= 16'hFD50;    16'd36553: out <= 16'hFC9D;    16'd36554: out <= 16'hFD0F;    16'd36555: out <= 16'h02BB;
    16'd36556: out <= 16'h019F;    16'd36557: out <= 16'h0380;    16'd36558: out <= 16'h049E;    16'd36559: out <= 16'h0A08;
    16'd36560: out <= 16'h0A00;    16'd36561: out <= 16'h0043;    16'd36562: out <= 16'h0338;    16'd36563: out <= 16'h0BD6;
    16'd36564: out <= 16'h0385;    16'd36565: out <= 16'h058E;    16'd36566: out <= 16'h041F;    16'd36567: out <= 16'h01FD;
    16'd36568: out <= 16'h050B;    16'd36569: out <= 16'h0273;    16'd36570: out <= 16'hF9D5;    16'd36571: out <= 16'h0347;
    16'd36572: out <= 16'h0764;    16'd36573: out <= 16'h0710;    16'd36574: out <= 16'h0243;    16'd36575: out <= 16'h0584;
    16'd36576: out <= 16'h02AA;    16'd36577: out <= 16'h078A;    16'd36578: out <= 16'h0153;    16'd36579: out <= 16'h099D;
    16'd36580: out <= 16'h088B;    16'd36581: out <= 16'h09BA;    16'd36582: out <= 16'h0618;    16'd36583: out <= 16'h0800;
    16'd36584: out <= 16'h0DDB;    16'd36585: out <= 16'h02D0;    16'd36586: out <= 16'h01DD;    16'd36587: out <= 16'hFACB;
    16'd36588: out <= 16'h00FB;    16'd36589: out <= 16'hF477;    16'd36590: out <= 16'h0154;    16'd36591: out <= 16'h0189;
    16'd36592: out <= 16'hFD5C;    16'd36593: out <= 16'hFD94;    16'd36594: out <= 16'hFF77;    16'd36595: out <= 16'hFE4B;
    16'd36596: out <= 16'h01E4;    16'd36597: out <= 16'hFD05;    16'd36598: out <= 16'h016D;    16'd36599: out <= 16'h0000;
    16'd36600: out <= 16'hFF4B;    16'd36601: out <= 16'hFEF9;    16'd36602: out <= 16'h00E7;    16'd36603: out <= 16'h00E8;
    16'd36604: out <= 16'hFD0E;    16'd36605: out <= 16'h043D;    16'd36606: out <= 16'h0587;    16'd36607: out <= 16'h0562;
    16'd36608: out <= 16'h016D;    16'd36609: out <= 16'hFE7F;    16'd36610: out <= 16'hFE9B;    16'd36611: out <= 16'hFB44;
    16'd36612: out <= 16'h013E;    16'd36613: out <= 16'h0148;    16'd36614: out <= 16'h0197;    16'd36615: out <= 16'h04EE;
    16'd36616: out <= 16'h0298;    16'd36617: out <= 16'h038C;    16'd36618: out <= 16'h03F8;    16'd36619: out <= 16'h01ED;
    16'd36620: out <= 16'h0159;    16'd36621: out <= 16'h0133;    16'd36622: out <= 16'hFD17;    16'd36623: out <= 16'h021E;
    16'd36624: out <= 16'hFD14;    16'd36625: out <= 16'h00A6;    16'd36626: out <= 16'h0141;    16'd36627: out <= 16'hFAB2;
    16'd36628: out <= 16'hFCDF;    16'd36629: out <= 16'h0167;    16'd36630: out <= 16'hFD21;    16'd36631: out <= 16'h007E;
    16'd36632: out <= 16'hFD62;    16'd36633: out <= 16'h0370;    16'd36634: out <= 16'h04C0;    16'd36635: out <= 16'h0DA6;
    16'd36636: out <= 16'h0390;    16'd36637: out <= 16'h0236;    16'd36638: out <= 16'h0514;    16'd36639: out <= 16'hFEB0;
    16'd36640: out <= 16'h07CB;    16'd36641: out <= 16'h0050;    16'd36642: out <= 16'hFE37;    16'd36643: out <= 16'h0E2C;
    16'd36644: out <= 16'h0014;    16'd36645: out <= 16'h04E7;    16'd36646: out <= 16'h01E5;    16'd36647: out <= 16'h0691;
    16'd36648: out <= 16'h05A9;    16'd36649: out <= 16'h073C;    16'd36650: out <= 16'h010B;    16'd36651: out <= 16'h04D2;
    16'd36652: out <= 16'h078E;    16'd36653: out <= 16'hFE4B;    16'd36654: out <= 16'hFFA1;    16'd36655: out <= 16'hFDB3;
    16'd36656: out <= 16'h0896;    16'd36657: out <= 16'h04E7;    16'd36658: out <= 16'h0385;    16'd36659: out <= 16'hFBD8;
    16'd36660: out <= 16'h06F5;    16'd36661: out <= 16'h0441;    16'd36662: out <= 16'h0034;    16'd36663: out <= 16'h05D0;
    16'd36664: out <= 16'h08A9;    16'd36665: out <= 16'h00BE;    16'd36666: out <= 16'h05CC;    16'd36667: out <= 16'h055A;
    16'd36668: out <= 16'h08C1;    16'd36669: out <= 16'h0470;    16'd36670: out <= 16'h03AC;    16'd36671: out <= 16'h0370;
    16'd36672: out <= 16'hFC28;    16'd36673: out <= 16'h0491;    16'd36674: out <= 16'h0375;    16'd36675: out <= 16'hFED5;
    16'd36676: out <= 16'h0337;    16'd36677: out <= 16'h020F;    16'd36678: out <= 16'h09DF;    16'd36679: out <= 16'h0307;
    16'd36680: out <= 16'h01D4;    16'd36681: out <= 16'hFE6B;    16'd36682: out <= 16'h0492;    16'd36683: out <= 16'h0632;
    16'd36684: out <= 16'h020B;    16'd36685: out <= 16'h0547;    16'd36686: out <= 16'h0044;    16'd36687: out <= 16'h03D9;
    16'd36688: out <= 16'h0180;    16'd36689: out <= 16'h0527;    16'd36690: out <= 16'h0123;    16'd36691: out <= 16'hFDC2;
    16'd36692: out <= 16'h01FE;    16'd36693: out <= 16'h0213;    16'd36694: out <= 16'h036D;    16'd36695: out <= 16'h0C3C;
    16'd36696: out <= 16'h0A3E;    16'd36697: out <= 16'h0398;    16'd36698: out <= 16'h01DD;    16'd36699: out <= 16'h07C4;
    16'd36700: out <= 16'h013D;    16'd36701: out <= 16'h0411;    16'd36702: out <= 16'h0460;    16'd36703: out <= 16'h02A9;
    16'd36704: out <= 16'h02CC;    16'd36705: out <= 16'h0C5B;    16'd36706: out <= 16'h0377;    16'd36707: out <= 16'h0324;
    16'd36708: out <= 16'h00FE;    16'd36709: out <= 16'hFFFA;    16'd36710: out <= 16'hFF49;    16'd36711: out <= 16'hF9CD;
    16'd36712: out <= 16'h0449;    16'd36713: out <= 16'hFC19;    16'd36714: out <= 16'h03F4;    16'd36715: out <= 16'hF928;
    16'd36716: out <= 16'h02F0;    16'd36717: out <= 16'h03B3;    16'd36718: out <= 16'h0360;    16'd36719: out <= 16'h09B8;
    16'd36720: out <= 16'h01F4;    16'd36721: out <= 16'h0254;    16'd36722: out <= 16'h02BF;    16'd36723: out <= 16'hFC1F;
    16'd36724: out <= 16'h00CD;    16'd36725: out <= 16'hFFD7;    16'd36726: out <= 16'h0361;    16'd36727: out <= 16'hFF37;
    16'd36728: out <= 16'h09AC;    16'd36729: out <= 16'h0809;    16'd36730: out <= 16'h0928;    16'd36731: out <= 16'h03DC;
    16'd36732: out <= 16'h0A27;    16'd36733: out <= 16'h0A15;    16'd36734: out <= 16'h0942;    16'd36735: out <= 16'h00C7;
    16'd36736: out <= 16'h06F3;    16'd36737: out <= 16'h00A7;    16'd36738: out <= 16'h01DD;    16'd36739: out <= 16'h05A4;
    16'd36740: out <= 16'h0548;    16'd36741: out <= 16'hFE41;    16'd36742: out <= 16'h028A;    16'd36743: out <= 16'hFB90;
    16'd36744: out <= 16'h01F8;    16'd36745: out <= 16'h05BF;    16'd36746: out <= 16'h088F;    16'd36747: out <= 16'hFFC3;
    16'd36748: out <= 16'h0570;    16'd36749: out <= 16'h021A;    16'd36750: out <= 16'h028F;    16'd36751: out <= 16'h0528;
    16'd36752: out <= 16'hFF3C;    16'd36753: out <= 16'h00B9;    16'd36754: out <= 16'h03A8;    16'd36755: out <= 16'h00A4;
    16'd36756: out <= 16'h07F3;    16'd36757: out <= 16'h05AC;    16'd36758: out <= 16'h0377;    16'd36759: out <= 16'h05AF;
    16'd36760: out <= 16'h019F;    16'd36761: out <= 16'h05F4;    16'd36762: out <= 16'h02C1;    16'd36763: out <= 16'h0360;
    16'd36764: out <= 16'h06DC;    16'd36765: out <= 16'h0333;    16'd36766: out <= 16'h000B;    16'd36767: out <= 16'h0190;
    16'd36768: out <= 16'hFE33;    16'd36769: out <= 16'h03FE;    16'd36770: out <= 16'h03BD;    16'd36771: out <= 16'h0A48;
    16'd36772: out <= 16'h0AD5;    16'd36773: out <= 16'h005B;    16'd36774: out <= 16'h05C6;    16'd36775: out <= 16'h034F;
    16'd36776: out <= 16'h0366;    16'd36777: out <= 16'h0507;    16'd36778: out <= 16'h03C8;    16'd36779: out <= 16'hFB53;
    16'd36780: out <= 16'h0202;    16'd36781: out <= 16'h01C4;    16'd36782: out <= 16'h0449;    16'd36783: out <= 16'h03BF;
    16'd36784: out <= 16'hF913;    16'd36785: out <= 16'h091B;    16'd36786: out <= 16'h01DE;    16'd36787: out <= 16'h0434;
    16'd36788: out <= 16'h0A87;    16'd36789: out <= 16'h01D5;    16'd36790: out <= 16'h06D0;    16'd36791: out <= 16'hFD7F;
    16'd36792: out <= 16'h0AAA;    16'd36793: out <= 16'h061E;    16'd36794: out <= 16'h0CDA;    16'd36795: out <= 16'h03A3;
    16'd36796: out <= 16'h054A;    16'd36797: out <= 16'h06F0;    16'd36798: out <= 16'h01B8;    16'd36799: out <= 16'h066D;
    16'd36800: out <= 16'h053E;    16'd36801: out <= 16'hFDDE;    16'd36802: out <= 16'h075D;    16'd36803: out <= 16'h046F;
    16'd36804: out <= 16'hFF68;    16'd36805: out <= 16'h0758;    16'd36806: out <= 16'h05B9;    16'd36807: out <= 16'h08CF;
    16'd36808: out <= 16'h04A2;    16'd36809: out <= 16'h044A;    16'd36810: out <= 16'h032B;    16'd36811: out <= 16'hFE45;
    16'd36812: out <= 16'hFD47;    16'd36813: out <= 16'h003A;    16'd36814: out <= 16'h0762;    16'd36815: out <= 16'h03F1;
    16'd36816: out <= 16'h004D;    16'd36817: out <= 16'h0926;    16'd36818: out <= 16'h04ED;    16'd36819: out <= 16'h04FA;
    16'd36820: out <= 16'h0779;    16'd36821: out <= 16'h0ABA;    16'd36822: out <= 16'h0585;    16'd36823: out <= 16'h01DD;
    16'd36824: out <= 16'h009D;    16'd36825: out <= 16'h00F0;    16'd36826: out <= 16'hFF39;    16'd36827: out <= 16'h004A;
    16'd36828: out <= 16'h03FA;    16'd36829: out <= 16'hFF8F;    16'd36830: out <= 16'h0640;    16'd36831: out <= 16'h045E;
    16'd36832: out <= 16'h0174;    16'd36833: out <= 16'h017D;    16'd36834: out <= 16'h03C7;    16'd36835: out <= 16'hFFB0;
    16'd36836: out <= 16'h0600;    16'd36837: out <= 16'h0424;    16'd36838: out <= 16'h0903;    16'd36839: out <= 16'h0785;
    16'd36840: out <= 16'h067F;    16'd36841: out <= 16'h01B8;    16'd36842: out <= 16'h0696;    16'd36843: out <= 16'hFFF1;
    16'd36844: out <= 16'hFE13;    16'd36845: out <= 16'h015A;    16'd36846: out <= 16'hFFFE;    16'd36847: out <= 16'hFE1C;
    16'd36848: out <= 16'h04D6;    16'd36849: out <= 16'h06E0;    16'd36850: out <= 16'h030E;    16'd36851: out <= 16'hFAE9;
    16'd36852: out <= 16'hFE43;    16'd36853: out <= 16'h00C1;    16'd36854: out <= 16'hFCA2;    16'd36855: out <= 16'h005F;
    16'd36856: out <= 16'h0821;    16'd36857: out <= 16'h0269;    16'd36858: out <= 16'hFF4D;    16'd36859: out <= 16'h0374;
    16'd36860: out <= 16'h04B2;    16'd36861: out <= 16'hFF01;    16'd36862: out <= 16'hFB16;    16'd36863: out <= 16'hFD8B;
    16'd36864: out <= 16'h001C;    16'd36865: out <= 16'hFF93;    16'd36866: out <= 16'hFB4E;    16'd36867: out <= 16'hFAD8;
    16'd36868: out <= 16'h035E;    16'd36869: out <= 16'h0571;    16'd36870: out <= 16'h04CB;    16'd36871: out <= 16'hFDE9;
    16'd36872: out <= 16'h0400;    16'd36873: out <= 16'hFCDF;    16'd36874: out <= 16'h02B9;    16'd36875: out <= 16'h03B3;
    16'd36876: out <= 16'hFC97;    16'd36877: out <= 16'h0262;    16'd36878: out <= 16'h02E3;    16'd36879: out <= 16'hFD5C;
    16'd36880: out <= 16'h020C;    16'd36881: out <= 16'hFC94;    16'd36882: out <= 16'h0369;    16'd36883: out <= 16'hFCCC;
    16'd36884: out <= 16'h0258;    16'd36885: out <= 16'hFE7A;    16'd36886: out <= 16'hFC53;    16'd36887: out <= 16'hFE0A;
    16'd36888: out <= 16'h028C;    16'd36889: out <= 16'h0482;    16'd36890: out <= 16'h01F4;    16'd36891: out <= 16'h033C;
    16'd36892: out <= 16'h047B;    16'd36893: out <= 16'h0642;    16'd36894: out <= 16'h090C;    16'd36895: out <= 16'hFF7D;
    16'd36896: out <= 16'h04EF;    16'd36897: out <= 16'h0301;    16'd36898: out <= 16'h0952;    16'd36899: out <= 16'hFFE8;
    16'd36900: out <= 16'h050C;    16'd36901: out <= 16'h0515;    16'd36902: out <= 16'h0459;    16'd36903: out <= 16'h03F5;
    16'd36904: out <= 16'h0577;    16'd36905: out <= 16'h0947;    16'd36906: out <= 16'h0670;    16'd36907: out <= 16'h03B8;
    16'd36908: out <= 16'h065A;    16'd36909: out <= 16'h061C;    16'd36910: out <= 16'h02DA;    16'd36911: out <= 16'hFF27;
    16'd36912: out <= 16'h0677;    16'd36913: out <= 16'h04E0;    16'd36914: out <= 16'h0982;    16'd36915: out <= 16'hFFCF;
    16'd36916: out <= 16'h02EA;    16'd36917: out <= 16'h0586;    16'd36918: out <= 16'h0794;    16'd36919: out <= 16'h0C05;
    16'd36920: out <= 16'h02ED;    16'd36921: out <= 16'h04AB;    16'd36922: out <= 16'h04A8;    16'd36923: out <= 16'hFB26;
    16'd36924: out <= 16'h02A2;    16'd36925: out <= 16'hFE18;    16'd36926: out <= 16'hFE79;    16'd36927: out <= 16'hFF3E;
    16'd36928: out <= 16'h0433;    16'd36929: out <= 16'h0144;    16'd36930: out <= 16'h0814;    16'd36931: out <= 16'h06B2;
    16'd36932: out <= 16'h089F;    16'd36933: out <= 16'h00A3;    16'd36934: out <= 16'h028F;    16'd36935: out <= 16'h02FC;
    16'd36936: out <= 16'h0210;    16'd36937: out <= 16'hFDB0;    16'd36938: out <= 16'h017C;    16'd36939: out <= 16'h0426;
    16'd36940: out <= 16'h0716;    16'd36941: out <= 16'h03E8;    16'd36942: out <= 16'h0061;    16'd36943: out <= 16'h053B;
    16'd36944: out <= 16'h0648;    16'd36945: out <= 16'h051A;    16'd36946: out <= 16'h04C2;    16'd36947: out <= 16'h005C;
    16'd36948: out <= 16'h0644;    16'd36949: out <= 16'h0D96;    16'd36950: out <= 16'h0202;    16'd36951: out <= 16'h059C;
    16'd36952: out <= 16'h0219;    16'd36953: out <= 16'hFEAC;    16'd36954: out <= 16'h0229;    16'd36955: out <= 16'h03DB;
    16'd36956: out <= 16'h02B4;    16'd36957: out <= 16'h0494;    16'd36958: out <= 16'h05B1;    16'd36959: out <= 16'hF98F;
    16'd36960: out <= 16'h022A;    16'd36961: out <= 16'h0284;    16'd36962: out <= 16'h0944;    16'd36963: out <= 16'hFDD1;
    16'd36964: out <= 16'h072C;    16'd36965: out <= 16'h035D;    16'd36966: out <= 16'h0278;    16'd36967: out <= 16'h07BF;
    16'd36968: out <= 16'h057E;    16'd36969: out <= 16'hFB3F;    16'd36970: out <= 16'h095E;    16'd36971: out <= 16'hFEEE;
    16'd36972: out <= 16'h00CF;    16'd36973: out <= 16'h01F0;    16'd36974: out <= 16'hFFF5;    16'd36975: out <= 16'h049A;
    16'd36976: out <= 16'h036C;    16'd36977: out <= 16'h05F8;    16'd36978: out <= 16'hFD8C;    16'd36979: out <= 16'h02F9;
    16'd36980: out <= 16'h0341;    16'd36981: out <= 16'hFE96;    16'd36982: out <= 16'hFF3D;    16'd36983: out <= 16'h017A;
    16'd36984: out <= 16'h0501;    16'd36985: out <= 16'h052E;    16'd36986: out <= 16'h05CA;    16'd36987: out <= 16'h053F;
    16'd36988: out <= 16'h00DF;    16'd36989: out <= 16'h0318;    16'd36990: out <= 16'h06D4;    16'd36991: out <= 16'hF839;
    16'd36992: out <= 16'hFEFE;    16'd36993: out <= 16'h01E2;    16'd36994: out <= 16'hFF1F;    16'd36995: out <= 16'hFFEC;
    16'd36996: out <= 16'h0286;    16'd36997: out <= 16'h00DC;    16'd36998: out <= 16'hFCAA;    16'd36999: out <= 16'hFF15;
    16'd37000: out <= 16'h05B8;    16'd37001: out <= 16'h03E3;    16'd37002: out <= 16'h01D2;    16'd37003: out <= 16'hFD43;
    16'd37004: out <= 16'hFC5E;    16'd37005: out <= 16'h0266;    16'd37006: out <= 16'h0663;    16'd37007: out <= 16'h0999;
    16'd37008: out <= 16'h06A7;    16'd37009: out <= 16'h0941;    16'd37010: out <= 16'hFFE6;    16'd37011: out <= 16'hFF78;
    16'd37012: out <= 16'hFE45;    16'd37013: out <= 16'h0768;    16'd37014: out <= 16'h0514;    16'd37015: out <= 16'h0447;
    16'd37016: out <= 16'h0042;    16'd37017: out <= 16'hFF60;    16'd37018: out <= 16'h0492;    16'd37019: out <= 16'h06B6;
    16'd37020: out <= 16'h0A1B;    16'd37021: out <= 16'hFC24;    16'd37022: out <= 16'h069F;    16'd37023: out <= 16'h070B;
    16'd37024: out <= 16'h046D;    16'd37025: out <= 16'h0625;    16'd37026: out <= 16'h0807;    16'd37027: out <= 16'hFF44;
    16'd37028: out <= 16'h03B9;    16'd37029: out <= 16'h05C6;    16'd37030: out <= 16'h0474;    16'd37031: out <= 16'h0334;
    16'd37032: out <= 16'h0485;    16'd37033: out <= 16'h0175;    16'd37034: out <= 16'h02B2;    16'd37035: out <= 16'h02D8;
    16'd37036: out <= 16'hFEAB;    16'd37037: out <= 16'h0522;    16'd37038: out <= 16'h05C5;    16'd37039: out <= 16'hFF0D;
    16'd37040: out <= 16'h0510;    16'd37041: out <= 16'h0140;    16'd37042: out <= 16'h092B;    16'd37043: out <= 16'h0ED3;
    16'd37044: out <= 16'h06F3;    16'd37045: out <= 16'h0300;    16'd37046: out <= 16'h04E9;    16'd37047: out <= 16'h0D79;
    16'd37048: out <= 16'h04E9;    16'd37049: out <= 16'h0642;    16'd37050: out <= 16'h0728;    16'd37051: out <= 16'h0B05;
    16'd37052: out <= 16'hFBEE;    16'd37053: out <= 16'h03DE;    16'd37054: out <= 16'h02D0;    16'd37055: out <= 16'h0478;
    16'd37056: out <= 16'h08BD;    16'd37057: out <= 16'h06FC;    16'd37058: out <= 16'hFDE3;    16'd37059: out <= 16'h055D;
    16'd37060: out <= 16'h06B0;    16'd37061: out <= 16'h0293;    16'd37062: out <= 16'hFF54;    16'd37063: out <= 16'h0176;
    16'd37064: out <= 16'h07F1;    16'd37065: out <= 16'h025E;    16'd37066: out <= 16'h0778;    16'd37067: out <= 16'h03EF;
    16'd37068: out <= 16'h05EB;    16'd37069: out <= 16'hFE63;    16'd37070: out <= 16'hF948;    16'd37071: out <= 16'h043B;
    16'd37072: out <= 16'hFE82;    16'd37073: out <= 16'h052E;    16'd37074: out <= 16'h00A1;    16'd37075: out <= 16'h020D;
    16'd37076: out <= 16'h02E4;    16'd37077: out <= 16'h0903;    16'd37078: out <= 16'h002C;    16'd37079: out <= 16'h00E2;
    16'd37080: out <= 16'h03D4;    16'd37081: out <= 16'h013A;    16'd37082: out <= 16'hFB92;    16'd37083: out <= 16'hF99E;
    16'd37084: out <= 16'h06AD;    16'd37085: out <= 16'h02B2;    16'd37086: out <= 16'hFE6B;    16'd37087: out <= 16'h07FA;
    16'd37088: out <= 16'h006E;    16'd37089: out <= 16'h0A3E;    16'd37090: out <= 16'h04AF;    16'd37091: out <= 16'h057C;
    16'd37092: out <= 16'h0186;    16'd37093: out <= 16'h030A;    16'd37094: out <= 16'h0023;    16'd37095: out <= 16'h065A;
    16'd37096: out <= 16'hFC3C;    16'd37097: out <= 16'h06BF;    16'd37098: out <= 16'h00D0;    16'd37099: out <= 16'h00F2;
    16'd37100: out <= 16'hFD45;    16'd37101: out <= 16'hFBEB;    16'd37102: out <= 16'hFE4F;    16'd37103: out <= 16'h0150;
    16'd37104: out <= 16'hF9FA;    16'd37105: out <= 16'h00CE;    16'd37106: out <= 16'hFBC5;    16'd37107: out <= 16'h0108;
    16'd37108: out <= 16'h05A8;    16'd37109: out <= 16'hFCAE;    16'd37110: out <= 16'hFF78;    16'd37111: out <= 16'hFCA3;
    16'd37112: out <= 16'h051B;    16'd37113: out <= 16'hFE6C;    16'd37114: out <= 16'hFD73;    16'd37115: out <= 16'hFF96;
    16'd37116: out <= 16'hFDBD;    16'd37117: out <= 16'hFDC4;    16'd37118: out <= 16'hFC1B;    16'd37119: out <= 16'h069F;
    16'd37120: out <= 16'hFB04;    16'd37121: out <= 16'hFD42;    16'd37122: out <= 16'h0173;    16'd37123: out <= 16'hFF18;
    16'd37124: out <= 16'h030A;    16'd37125: out <= 16'hF68D;    16'd37126: out <= 16'hFD17;    16'd37127: out <= 16'hF3D7;
    16'd37128: out <= 16'hFE29;    16'd37129: out <= 16'hFD04;    16'd37130: out <= 16'hFF67;    16'd37131: out <= 16'h000A;
    16'd37132: out <= 16'hF694;    16'd37133: out <= 16'h01EA;    16'd37134: out <= 16'h06AC;    16'd37135: out <= 16'hFF66;
    16'd37136: out <= 16'hFE9A;    16'd37137: out <= 16'hFF7C;    16'd37138: out <= 16'h01CB;    16'd37139: out <= 16'hF8E0;
    16'd37140: out <= 16'h029B;    16'd37141: out <= 16'h0377;    16'd37142: out <= 16'hFE4C;    16'd37143: out <= 16'hFC0B;
    16'd37144: out <= 16'h03A0;    16'd37145: out <= 16'hFEB0;    16'd37146: out <= 16'h0469;    16'd37147: out <= 16'h0297;
    16'd37148: out <= 16'h034B;    16'd37149: out <= 16'h0784;    16'd37150: out <= 16'h0925;    16'd37151: out <= 16'hFF67;
    16'd37152: out <= 16'h0427;    16'd37153: out <= 16'h05D5;    16'd37154: out <= 16'h0547;    16'd37155: out <= 16'hFEDE;
    16'd37156: out <= 16'h09FD;    16'd37157: out <= 16'h0552;    16'd37158: out <= 16'h01FD;    16'd37159: out <= 16'h0AAF;
    16'd37160: out <= 16'hFF42;    16'd37161: out <= 16'h0564;    16'd37162: out <= 16'h0047;    16'd37163: out <= 16'h0483;
    16'd37164: out <= 16'h09C6;    16'd37165: out <= 16'h07BB;    16'd37166: out <= 16'h01B4;    16'd37167: out <= 16'h0298;
    16'd37168: out <= 16'h02EA;    16'd37169: out <= 16'h0806;    16'd37170: out <= 16'h0408;    16'd37171: out <= 16'h0232;
    16'd37172: out <= 16'h0B42;    16'd37173: out <= 16'h028F;    16'd37174: out <= 16'h063C;    16'd37175: out <= 16'h08B2;
    16'd37176: out <= 16'hFDFA;    16'd37177: out <= 16'hF5F5;    16'd37178: out <= 16'h056D;    16'd37179: out <= 16'h0078;
    16'd37180: out <= 16'hFF8E;    16'd37181: out <= 16'h06D0;    16'd37182: out <= 16'h0020;    16'd37183: out <= 16'h0636;
    16'd37184: out <= 16'h0775;    16'd37185: out <= 16'h0675;    16'd37186: out <= 16'h0A92;    16'd37187: out <= 16'h0366;
    16'd37188: out <= 16'h07C8;    16'd37189: out <= 16'h0387;    16'd37190: out <= 16'h050D;    16'd37191: out <= 16'h0837;
    16'd37192: out <= 16'h0250;    16'd37193: out <= 16'h0DA1;    16'd37194: out <= 16'h0278;    16'd37195: out <= 16'hFB8E;
    16'd37196: out <= 16'hFE84;    16'd37197: out <= 16'h06A3;    16'd37198: out <= 16'h06D0;    16'd37199: out <= 16'h027B;
    16'd37200: out <= 16'h05FF;    16'd37201: out <= 16'hFFBC;    16'd37202: out <= 16'h02FA;    16'd37203: out <= 16'h078F;
    16'd37204: out <= 16'h064A;    16'd37205: out <= 16'h0961;    16'd37206: out <= 16'h0738;    16'd37207: out <= 16'hFD5B;
    16'd37208: out <= 16'h0020;    16'd37209: out <= 16'h0548;    16'd37210: out <= 16'hFC75;    16'd37211: out <= 16'h0B60;
    16'd37212: out <= 16'h04C3;    16'd37213: out <= 16'h0445;    16'd37214: out <= 16'h0D53;    16'd37215: out <= 16'hFDD5;
    16'd37216: out <= 16'hFC1D;    16'd37217: out <= 16'h0846;    16'd37218: out <= 16'h02DF;    16'd37219: out <= 16'h03B2;
    16'd37220: out <= 16'h002E;    16'd37221: out <= 16'h0028;    16'd37222: out <= 16'h0386;    16'd37223: out <= 16'hFEF1;
    16'd37224: out <= 16'h0130;    16'd37225: out <= 16'hF889;    16'd37226: out <= 16'hFA85;    16'd37227: out <= 16'hF5C2;
    16'd37228: out <= 16'h0511;    16'd37229: out <= 16'h0133;    16'd37230: out <= 16'h068F;    16'd37231: out <= 16'h067C;
    16'd37232: out <= 16'h03B0;    16'd37233: out <= 16'h00BE;    16'd37234: out <= 16'h029E;    16'd37235: out <= 16'h03E5;
    16'd37236: out <= 16'hFC64;    16'd37237: out <= 16'hFE61;    16'd37238: out <= 16'h01FE;    16'd37239: out <= 16'h04F4;
    16'd37240: out <= 16'hFDF6;    16'd37241: out <= 16'h0975;    16'd37242: out <= 16'h0777;    16'd37243: out <= 16'h0731;
    16'd37244: out <= 16'hFF99;    16'd37245: out <= 16'hFFD7;    16'd37246: out <= 16'h0206;    16'd37247: out <= 16'h01D3;
    16'd37248: out <= 16'h00E2;    16'd37249: out <= 16'hF8F6;    16'd37250: out <= 16'hFD7B;    16'd37251: out <= 16'hFBE7;
    16'd37252: out <= 16'h0314;    16'd37253: out <= 16'h013D;    16'd37254: out <= 16'hFD21;    16'd37255: out <= 16'hFD5C;
    16'd37256: out <= 16'h03A7;    16'd37257: out <= 16'hFF83;    16'd37258: out <= 16'h035E;    16'd37259: out <= 16'h02F0;
    16'd37260: out <= 16'h0119;    16'd37261: out <= 16'h02EB;    16'd37262: out <= 16'h0789;    16'd37263: out <= 16'h02A3;
    16'd37264: out <= 16'hFC7F;    16'd37265: out <= 16'h0267;    16'd37266: out <= 16'hFC9C;    16'd37267: out <= 16'hFCE1;
    16'd37268: out <= 16'h03D8;    16'd37269: out <= 16'h02CA;    16'd37270: out <= 16'hFF81;    16'd37271: out <= 16'h00E4;
    16'd37272: out <= 16'h0437;    16'd37273: out <= 16'h0708;    16'd37274: out <= 16'hFCA5;    16'd37275: out <= 16'h09F5;
    16'd37276: out <= 16'h0493;    16'd37277: out <= 16'h0201;    16'd37278: out <= 16'h053C;    16'd37279: out <= 16'h0510;
    16'd37280: out <= 16'hFD11;    16'd37281: out <= 16'h04F3;    16'd37282: out <= 16'h0259;    16'd37283: out <= 16'h0D88;
    16'd37284: out <= 16'h0328;    16'd37285: out <= 16'hFF58;    16'd37286: out <= 16'h0B50;    16'd37287: out <= 16'h0574;
    16'd37288: out <= 16'h0CF7;    16'd37289: out <= 16'h02E4;    16'd37290: out <= 16'h00D9;    16'd37291: out <= 16'h0464;
    16'd37292: out <= 16'h05D0;    16'd37293: out <= 16'hFFCF;    16'd37294: out <= 16'h06EE;    16'd37295: out <= 16'hF90F;
    16'd37296: out <= 16'h0779;    16'd37297: out <= 16'h07AF;    16'd37298: out <= 16'h05BE;    16'd37299: out <= 16'h0906;
    16'd37300: out <= 16'h0A83;    16'd37301: out <= 16'h02D5;    16'd37302: out <= 16'h0496;    16'd37303: out <= 16'h0C5B;
    16'd37304: out <= 16'h0575;    16'd37305: out <= 16'h05F9;    16'd37306: out <= 16'h0146;    16'd37307: out <= 16'h063A;
    16'd37308: out <= 16'h0162;    16'd37309: out <= 16'h03E9;    16'd37310: out <= 16'h00B6;    16'd37311: out <= 16'h02FF;
    16'd37312: out <= 16'h07AD;    16'd37313: out <= 16'h0154;    16'd37314: out <= 16'h000F;    16'd37315: out <= 16'h0882;
    16'd37316: out <= 16'h062E;    16'd37317: out <= 16'h0066;    16'd37318: out <= 16'h010A;    16'd37319: out <= 16'h057B;
    16'd37320: out <= 16'h070C;    16'd37321: out <= 16'h09C9;    16'd37322: out <= 16'h0B5B;    16'd37323: out <= 16'h06EC;
    16'd37324: out <= 16'h07FB;    16'd37325: out <= 16'h09AC;    16'd37326: out <= 16'h03A9;    16'd37327: out <= 16'h049E;
    16'd37328: out <= 16'h0735;    16'd37329: out <= 16'h06E2;    16'd37330: out <= 16'h04C0;    16'd37331: out <= 16'h0362;
    16'd37332: out <= 16'h01CF;    16'd37333: out <= 16'h0526;    16'd37334: out <= 16'h061A;    16'd37335: out <= 16'hFC8E;
    16'd37336: out <= 16'h059A;    16'd37337: out <= 16'hFE0C;    16'd37338: out <= 16'h01D7;    16'd37339: out <= 16'h023A;
    16'd37340: out <= 16'h029D;    16'd37341: out <= 16'h0268;    16'd37342: out <= 16'h03C1;    16'd37343: out <= 16'h02F1;
    16'd37344: out <= 16'h0572;    16'd37345: out <= 16'h014A;    16'd37346: out <= 16'h05D6;    16'd37347: out <= 16'h090E;
    16'd37348: out <= 16'h01B7;    16'd37349: out <= 16'h06CF;    16'd37350: out <= 16'h01CD;    16'd37351: out <= 16'h0451;
    16'd37352: out <= 16'hFE70;    16'd37353: out <= 16'hFC05;    16'd37354: out <= 16'hF671;    16'd37355: out <= 16'hFDE2;
    16'd37356: out <= 16'hFED2;    16'd37357: out <= 16'hFBA5;    16'd37358: out <= 16'hFF00;    16'd37359: out <= 16'h0223;
    16'd37360: out <= 16'hFA7D;    16'd37361: out <= 16'h0589;    16'd37362: out <= 16'hFA7A;    16'd37363: out <= 16'h00FB;
    16'd37364: out <= 16'hFDD6;    16'd37365: out <= 16'h0117;    16'd37366: out <= 16'h0219;    16'd37367: out <= 16'h027B;
    16'd37368: out <= 16'h04A0;    16'd37369: out <= 16'hFF07;    16'd37370: out <= 16'hFC05;    16'd37371: out <= 16'h009F;
    16'd37372: out <= 16'h00B8;    16'd37373: out <= 16'hFFCD;    16'd37374: out <= 16'hF99E;    16'd37375: out <= 16'h032D;
    16'd37376: out <= 16'h00B2;    16'd37377: out <= 16'h007B;    16'd37378: out <= 16'h006E;    16'd37379: out <= 16'h0331;
    16'd37380: out <= 16'h028B;    16'd37381: out <= 16'hFBA1;    16'd37382: out <= 16'hFEA7;    16'd37383: out <= 16'h067F;
    16'd37384: out <= 16'h03BD;    16'd37385: out <= 16'hFBA8;    16'd37386: out <= 16'hFDA6;    16'd37387: out <= 16'hFF01;
    16'd37388: out <= 16'hF9D1;    16'd37389: out <= 16'h0197;    16'd37390: out <= 16'h0348;    16'd37391: out <= 16'h03A4;
    16'd37392: out <= 16'h075D;    16'd37393: out <= 16'h022F;    16'd37394: out <= 16'h0078;    16'd37395: out <= 16'h0588;
    16'd37396: out <= 16'h003D;    16'd37397: out <= 16'h0123;    16'd37398: out <= 16'hFD00;    16'd37399: out <= 16'hFF5E;
    16'd37400: out <= 16'hFAE2;    16'd37401: out <= 16'hFF19;    16'd37402: out <= 16'h0173;    16'd37403: out <= 16'h04E0;
    16'd37404: out <= 16'h044A;    16'd37405: out <= 16'h03F4;    16'd37406: out <= 16'hFEEE;    16'd37407: out <= 16'h00E2;
    16'd37408: out <= 16'h04E0;    16'd37409: out <= 16'h01E3;    16'd37410: out <= 16'h00C6;    16'd37411: out <= 16'h03E5;
    16'd37412: out <= 16'h0491;    16'd37413: out <= 16'h06EC;    16'd37414: out <= 16'h0690;    16'd37415: out <= 16'h014F;
    16'd37416: out <= 16'h00D1;    16'd37417: out <= 16'h0752;    16'd37418: out <= 16'h0581;    16'd37419: out <= 16'hFD83;
    16'd37420: out <= 16'h03EF;    16'd37421: out <= 16'h0413;    16'd37422: out <= 16'h0436;    16'd37423: out <= 16'h0759;
    16'd37424: out <= 16'h0372;    16'd37425: out <= 16'hFFED;    16'd37426: out <= 16'h05E7;    16'd37427: out <= 16'hFD5B;
    16'd37428: out <= 16'h0265;    16'd37429: out <= 16'h0254;    16'd37430: out <= 16'h000B;    16'd37431: out <= 16'h0694;
    16'd37432: out <= 16'h0334;    16'd37433: out <= 16'h0435;    16'd37434: out <= 16'h07B8;    16'd37435: out <= 16'h0B19;
    16'd37436: out <= 16'h0290;    16'd37437: out <= 16'h079A;    16'd37438: out <= 16'h00D8;    16'd37439: out <= 16'h016B;
    16'd37440: out <= 16'h0034;    16'd37441: out <= 16'h03B0;    16'd37442: out <= 16'h06E3;    16'd37443: out <= 16'h01E1;
    16'd37444: out <= 16'h0595;    16'd37445: out <= 16'h07AD;    16'd37446: out <= 16'h0461;    16'd37447: out <= 16'h07E8;
    16'd37448: out <= 16'h03A6;    16'd37449: out <= 16'h0031;    16'd37450: out <= 16'h06A9;    16'd37451: out <= 16'h0721;
    16'd37452: out <= 16'h0487;    16'd37453: out <= 16'h05AA;    16'd37454: out <= 16'h0A2C;    16'd37455: out <= 16'h070B;
    16'd37456: out <= 16'h081B;    16'd37457: out <= 16'h026A;    16'd37458: out <= 16'h0546;    16'd37459: out <= 16'hFD22;
    16'd37460: out <= 16'h05C1;    16'd37461: out <= 16'h02DF;    16'd37462: out <= 16'hFDAC;    16'd37463: out <= 16'h05C4;
    16'd37464: out <= 16'h03B9;    16'd37465: out <= 16'h0067;    16'd37466: out <= 16'h07C6;    16'd37467: out <= 16'h00F0;
    16'd37468: out <= 16'h0179;    16'd37469: out <= 16'h0613;    16'd37470: out <= 16'h07EC;    16'd37471: out <= 16'hFD3B;
    16'd37472: out <= 16'hFEEA;    16'd37473: out <= 16'h0A52;    16'd37474: out <= 16'h06E6;    16'd37475: out <= 16'h0769;
    16'd37476: out <= 16'h0B8A;    16'd37477: out <= 16'h039B;    16'd37478: out <= 16'hFFEC;    16'd37479: out <= 16'hFD70;
    16'd37480: out <= 16'hFD8B;    16'd37481: out <= 16'h0415;    16'd37482: out <= 16'h0173;    16'd37483: out <= 16'h004C;
    16'd37484: out <= 16'h03C4;    16'd37485: out <= 16'h0210;    16'd37486: out <= 16'h04DB;    16'd37487: out <= 16'h078E;
    16'd37488: out <= 16'hFD7F;    16'd37489: out <= 16'h08A8;    16'd37490: out <= 16'h05D1;    16'd37491: out <= 16'h01FB;
    16'd37492: out <= 16'h001C;    16'd37493: out <= 16'h079C;    16'd37494: out <= 16'hF8FA;    16'd37495: out <= 16'h013B;
    16'd37496: out <= 16'h0089;    16'd37497: out <= 16'h00C7;    16'd37498: out <= 16'h019C;    16'd37499: out <= 16'h033E;
    16'd37500: out <= 16'h07A2;    16'd37501: out <= 16'h0111;    16'd37502: out <= 16'h03B3;    16'd37503: out <= 16'hFF29;
    16'd37504: out <= 16'hFF98;    16'd37505: out <= 16'hFA3A;    16'd37506: out <= 16'h0549;    16'd37507: out <= 16'h001B;
    16'd37508: out <= 16'hFA20;    16'd37509: out <= 16'h003F;    16'd37510: out <= 16'h037B;    16'd37511: out <= 16'h047A;
    16'd37512: out <= 16'hFCCD;    16'd37513: out <= 16'hFE42;    16'd37514: out <= 16'h0A06;    16'd37515: out <= 16'h0585;
    16'd37516: out <= 16'h0388;    16'd37517: out <= 16'h08F8;    16'd37518: out <= 16'h0239;    16'd37519: out <= 16'h0B28;
    16'd37520: out <= 16'h02B7;    16'd37521: out <= 16'h06F8;    16'd37522: out <= 16'h0264;    16'd37523: out <= 16'h0593;
    16'd37524: out <= 16'h03E2;    16'd37525: out <= 16'h036B;    16'd37526: out <= 16'h0498;    16'd37527: out <= 16'h0504;
    16'd37528: out <= 16'h08FC;    16'd37529: out <= 16'h0590;    16'd37530: out <= 16'h0750;    16'd37531: out <= 16'hFF13;
    16'd37532: out <= 16'h026D;    16'd37533: out <= 16'h01C9;    16'd37534: out <= 16'h04E9;    16'd37535: out <= 16'h0549;
    16'd37536: out <= 16'h0911;    16'd37537: out <= 16'h0B08;    16'd37538: out <= 16'h0261;    16'd37539: out <= 16'h04A5;
    16'd37540: out <= 16'hFD69;    16'd37541: out <= 16'hFD6C;    16'd37542: out <= 16'h032A;    16'd37543: out <= 16'h04B8;
    16'd37544: out <= 16'h0787;    16'd37545: out <= 16'h027B;    16'd37546: out <= 16'hFFB9;    16'd37547: out <= 16'h0657;
    16'd37548: out <= 16'h0684;    16'd37549: out <= 16'h05A3;    16'd37550: out <= 16'h03D0;    16'd37551: out <= 16'h01C9;
    16'd37552: out <= 16'h06CE;    16'd37553: out <= 16'h06AA;    16'd37554: out <= 16'h0014;    16'd37555: out <= 16'h0613;
    16'd37556: out <= 16'h05DC;    16'd37557: out <= 16'h04A5;    16'd37558: out <= 16'h07D8;    16'd37559: out <= 16'h0919;
    16'd37560: out <= 16'h09B7;    16'd37561: out <= 16'h0341;    16'd37562: out <= 16'h0B41;    16'd37563: out <= 16'h05BE;
    16'd37564: out <= 16'hFFCB;    16'd37565: out <= 16'hFE1D;    16'd37566: out <= 16'h0738;    16'd37567: out <= 16'h055C;
    16'd37568: out <= 16'h06A6;    16'd37569: out <= 16'h00A8;    16'd37570: out <= 16'h0377;    16'd37571: out <= 16'hFEEC;
    16'd37572: out <= 16'h0379;    16'd37573: out <= 16'h07A8;    16'd37574: out <= 16'hFFFC;    16'd37575: out <= 16'h062E;
    16'd37576: out <= 16'hFF45;    16'd37577: out <= 16'h0A8A;    16'd37578: out <= 16'h02D7;    16'd37579: out <= 16'h081B;
    16'd37580: out <= 16'h01A2;    16'd37581: out <= 16'h04C5;    16'd37582: out <= 16'h0156;    16'd37583: out <= 16'h0206;
    16'd37584: out <= 16'h08B2;    16'd37585: out <= 16'h070E;    16'd37586: out <= 16'hFFF3;    16'd37587: out <= 16'h0A0D;
    16'd37588: out <= 16'h057C;    16'd37589: out <= 16'h090B;    16'd37590: out <= 16'h0391;    16'd37591: out <= 16'hFCEE;
    16'd37592: out <= 16'hF86B;    16'd37593: out <= 16'hFD4D;    16'd37594: out <= 16'h010F;    16'd37595: out <= 16'h01EA;
    16'd37596: out <= 16'h004C;    16'd37597: out <= 16'h01B7;    16'd37598: out <= 16'hFFFD;    16'd37599: out <= 16'hFEE4;
    16'd37600: out <= 16'h042D;    16'd37601: out <= 16'h04E5;    16'd37602: out <= 16'h0B68;    16'd37603: out <= 16'h0423;
    16'd37604: out <= 16'h0159;    16'd37605: out <= 16'h027A;    16'd37606: out <= 16'h03E5;    16'd37607: out <= 16'h0114;
    16'd37608: out <= 16'h042D;    16'd37609: out <= 16'h00FE;    16'd37610: out <= 16'hFEB0;    16'd37611: out <= 16'h00A9;
    16'd37612: out <= 16'hFCEC;    16'd37613: out <= 16'h04FF;    16'd37614: out <= 16'hFA49;    16'd37615: out <= 16'h045E;
    16'd37616: out <= 16'hFCA5;    16'd37617: out <= 16'h03B9;    16'd37618: out <= 16'hFFA9;    16'd37619: out <= 16'h0097;
    16'd37620: out <= 16'hF835;    16'd37621: out <= 16'hFD11;    16'd37622: out <= 16'hFEFF;    16'd37623: out <= 16'h022C;
    16'd37624: out <= 16'hFBD4;    16'd37625: out <= 16'h04B9;    16'd37626: out <= 16'h027A;    16'd37627: out <= 16'hFA72;
    16'd37628: out <= 16'hFBAF;    16'd37629: out <= 16'h007C;    16'd37630: out <= 16'hFDC8;    16'd37631: out <= 16'hFED9;
    16'd37632: out <= 16'hFF43;    16'd37633: out <= 16'hFDBF;    16'd37634: out <= 16'hFF84;    16'd37635: out <= 16'h0141;
    16'd37636: out <= 16'h094C;    16'd37637: out <= 16'hFEB3;    16'd37638: out <= 16'hFEA6;    16'd37639: out <= 16'h0550;
    16'd37640: out <= 16'hFF13;    16'd37641: out <= 16'h00AF;    16'd37642: out <= 16'h01BC;    16'd37643: out <= 16'hFEEF;
    16'd37644: out <= 16'hFF2F;    16'd37645: out <= 16'h0051;    16'd37646: out <= 16'h0381;    16'd37647: out <= 16'hFE9D;
    16'd37648: out <= 16'h00D8;    16'd37649: out <= 16'h00BB;    16'd37650: out <= 16'hFC0C;    16'd37651: out <= 16'h0278;
    16'd37652: out <= 16'hF915;    16'd37653: out <= 16'h0069;    16'd37654: out <= 16'h00BE;    16'd37655: out <= 16'h01BD;
    16'd37656: out <= 16'hFD9B;    16'd37657: out <= 16'hFF02;    16'd37658: out <= 16'h05A1;    16'd37659: out <= 16'h0631;
    16'd37660: out <= 16'h087D;    16'd37661: out <= 16'h0675;    16'd37662: out <= 16'h04C3;    16'd37663: out <= 16'h0212;
    16'd37664: out <= 16'h0432;    16'd37665: out <= 16'h069E;    16'd37666: out <= 16'h0411;    16'd37667: out <= 16'h08AA;
    16'd37668: out <= 16'h0254;    16'd37669: out <= 16'h0959;    16'd37670: out <= 16'h0471;    16'd37671: out <= 16'hFE73;
    16'd37672: out <= 16'h0F22;    16'd37673: out <= 16'h0B67;    16'd37674: out <= 16'h0563;    16'd37675: out <= 16'h015E;
    16'd37676: out <= 16'h0016;    16'd37677: out <= 16'hFB7A;    16'd37678: out <= 16'h0C4A;    16'd37679: out <= 16'h0230;
    16'd37680: out <= 16'h0159;    16'd37681: out <= 16'h050A;    16'd37682: out <= 16'hF86D;    16'd37683: out <= 16'h02E0;
    16'd37684: out <= 16'h0151;    16'd37685: out <= 16'h03C2;    16'd37686: out <= 16'h065A;    16'd37687: out <= 16'h016A;
    16'd37688: out <= 16'h0202;    16'd37689: out <= 16'h06A0;    16'd37690: out <= 16'h0068;    16'd37691: out <= 16'h0656;
    16'd37692: out <= 16'h0B65;    16'd37693: out <= 16'hFFF1;    16'd37694: out <= 16'h008A;    16'd37695: out <= 16'h0633;
    16'd37696: out <= 16'h0529;    16'd37697: out <= 16'h00D2;    16'd37698: out <= 16'h07AD;    16'd37699: out <= 16'h0475;
    16'd37700: out <= 16'hFEE7;    16'd37701: out <= 16'h01A0;    16'd37702: out <= 16'h00B9;    16'd37703: out <= 16'h0381;
    16'd37704: out <= 16'h036D;    16'd37705: out <= 16'h07FA;    16'd37706: out <= 16'h0527;    16'd37707: out <= 16'h0645;
    16'd37708: out <= 16'h0392;    16'd37709: out <= 16'h0053;    16'd37710: out <= 16'h0881;    16'd37711: out <= 16'hFEA7;
    16'd37712: out <= 16'h09E1;    16'd37713: out <= 16'h04CC;    16'd37714: out <= 16'h005A;    16'd37715: out <= 16'h0597;
    16'd37716: out <= 16'h0436;    16'd37717: out <= 16'h01F6;    16'd37718: out <= 16'h032C;    16'd37719: out <= 16'h0910;
    16'd37720: out <= 16'h029D;    16'd37721: out <= 16'h000D;    16'd37722: out <= 16'h077A;    16'd37723: out <= 16'h0108;
    16'd37724: out <= 16'h0235;    16'd37725: out <= 16'h0B63;    16'd37726: out <= 16'h012B;    16'd37727: out <= 16'h0596;
    16'd37728: out <= 16'h007D;    16'd37729: out <= 16'h07EC;    16'd37730: out <= 16'h02E5;    16'd37731: out <= 16'h02F3;
    16'd37732: out <= 16'h0093;    16'd37733: out <= 16'hFD4E;    16'd37734: out <= 16'h036B;    16'd37735: out <= 16'h00FC;
    16'd37736: out <= 16'hFECB;    16'd37737: out <= 16'hFF9A;    16'd37738: out <= 16'h07C6;    16'd37739: out <= 16'h06E0;
    16'd37740: out <= 16'hFFF7;    16'd37741: out <= 16'h0359;    16'd37742: out <= 16'hFF57;    16'd37743: out <= 16'h08AF;
    16'd37744: out <= 16'h079A;    16'd37745: out <= 16'h07C8;    16'd37746: out <= 16'h0294;    16'd37747: out <= 16'h086E;
    16'd37748: out <= 16'hF9A0;    16'd37749: out <= 16'hFCFE;    16'd37750: out <= 16'hFF93;    16'd37751: out <= 16'h0020;
    16'd37752: out <= 16'hFEE2;    16'd37753: out <= 16'h0227;    16'd37754: out <= 16'h0C22;    16'd37755: out <= 16'h0321;
    16'd37756: out <= 16'h09DB;    16'd37757: out <= 16'h05B6;    16'd37758: out <= 16'h0227;    16'd37759: out <= 16'h055F;
    16'd37760: out <= 16'h037F;    16'd37761: out <= 16'h004C;    16'd37762: out <= 16'h0409;    16'd37763: out <= 16'hFEA0;
    16'd37764: out <= 16'hFCDE;    16'd37765: out <= 16'hFB5E;    16'd37766: out <= 16'h0654;    16'd37767: out <= 16'hFF87;
    16'd37768: out <= 16'h021D;    16'd37769: out <= 16'h017E;    16'd37770: out <= 16'hFC58;    16'd37771: out <= 16'hFEBD;
    16'd37772: out <= 16'h027E;    16'd37773: out <= 16'h0076;    16'd37774: out <= 16'h0CBE;    16'd37775: out <= 16'hFB6C;
    16'd37776: out <= 16'h0782;    16'd37777: out <= 16'h0332;    16'd37778: out <= 16'h0847;    16'd37779: out <= 16'h0308;
    16'd37780: out <= 16'h00FD;    16'd37781: out <= 16'h041B;    16'd37782: out <= 16'h03B4;    16'd37783: out <= 16'hFDC3;
    16'd37784: out <= 16'h0550;    16'd37785: out <= 16'hFF1C;    16'd37786: out <= 16'h0311;    16'd37787: out <= 16'h0265;
    16'd37788: out <= 16'h03A7;    16'd37789: out <= 16'h0822;    16'd37790: out <= 16'hFF32;    16'd37791: out <= 16'hFE28;
    16'd37792: out <= 16'h02F4;    16'd37793: out <= 16'h0964;    16'd37794: out <= 16'h049F;    16'd37795: out <= 16'h07D4;
    16'd37796: out <= 16'h0776;    16'd37797: out <= 16'h04F3;    16'd37798: out <= 16'h04A8;    16'd37799: out <= 16'h0843;
    16'd37800: out <= 16'h047F;    16'd37801: out <= 16'h0217;    16'd37802: out <= 16'hFCEC;    16'd37803: out <= 16'h09F5;
    16'd37804: out <= 16'h02D0;    16'd37805: out <= 16'h042D;    16'd37806: out <= 16'h07AD;    16'd37807: out <= 16'h00C9;
    16'd37808: out <= 16'h0500;    16'd37809: out <= 16'h0715;    16'd37810: out <= 16'h0301;    16'd37811: out <= 16'h01AE;
    16'd37812: out <= 16'h06DB;    16'd37813: out <= 16'h08AA;    16'd37814: out <= 16'h00CE;    16'd37815: out <= 16'h026E;
    16'd37816: out <= 16'h0289;    16'd37817: out <= 16'h03B9;    16'd37818: out <= 16'h0167;    16'd37819: out <= 16'h0642;
    16'd37820: out <= 16'h0484;    16'd37821: out <= 16'h0484;    16'd37822: out <= 16'h06C6;    16'd37823: out <= 16'h0877;
    16'd37824: out <= 16'h05BC;    16'd37825: out <= 16'hFF96;    16'd37826: out <= 16'h07D4;    16'd37827: out <= 16'h0930;
    16'd37828: out <= 16'h019B;    16'd37829: out <= 16'h0859;    16'd37830: out <= 16'h05F0;    16'd37831: out <= 16'h05D1;
    16'd37832: out <= 16'h0B70;    16'd37833: out <= 16'h0CF3;    16'd37834: out <= 16'h082F;    16'd37835: out <= 16'h014C;
    16'd37836: out <= 16'h0727;    16'd37837: out <= 16'h0119;    16'd37838: out <= 16'h027B;    16'd37839: out <= 16'h016C;
    16'd37840: out <= 16'h08A6;    16'd37841: out <= 16'hFC82;    16'd37842: out <= 16'h0275;    16'd37843: out <= 16'h0799;
    16'd37844: out <= 16'hFED5;    16'd37845: out <= 16'h040F;    16'd37846: out <= 16'h01EC;    16'd37847: out <= 16'h02A9;
    16'd37848: out <= 16'h06D0;    16'd37849: out <= 16'h0177;    16'd37850: out <= 16'h063F;    16'd37851: out <= 16'h037C;
    16'd37852: out <= 16'hFEE2;    16'd37853: out <= 16'h0105;    16'd37854: out <= 16'h01DF;    16'd37855: out <= 16'h0786;
    16'd37856: out <= 16'hFDFE;    16'd37857: out <= 16'h01F2;    16'd37858: out <= 16'h0129;    16'd37859: out <= 16'hFD9C;
    16'd37860: out <= 16'h073D;    16'd37861: out <= 16'h0B2A;    16'd37862: out <= 16'h0080;    16'd37863: out <= 16'h0241;
    16'd37864: out <= 16'hFF6F;    16'd37865: out <= 16'hFECB;    16'd37866: out <= 16'hFC80;    16'd37867: out <= 16'h02E7;
    16'd37868: out <= 16'hFDF5;    16'd37869: out <= 16'h0419;    16'd37870: out <= 16'h01E8;    16'd37871: out <= 16'h0297;
    16'd37872: out <= 16'hFDD3;    16'd37873: out <= 16'h01F0;    16'd37874: out <= 16'h00DB;    16'd37875: out <= 16'hFCF3;
    16'd37876: out <= 16'hFD51;    16'd37877: out <= 16'hFB76;    16'd37878: out <= 16'hFCB2;    16'd37879: out <= 16'h0438;
    16'd37880: out <= 16'h01DF;    16'd37881: out <= 16'hFF21;    16'd37882: out <= 16'h022E;    16'd37883: out <= 16'h0155;
    16'd37884: out <= 16'h05F1;    16'd37885: out <= 16'h0234;    16'd37886: out <= 16'hF009;    16'd37887: out <= 16'h01C6;
    16'd37888: out <= 16'h0106;    16'd37889: out <= 16'h015E;    16'd37890: out <= 16'h03C2;    16'd37891: out <= 16'h0404;
    16'd37892: out <= 16'h0070;    16'd37893: out <= 16'h015E;    16'd37894: out <= 16'h008E;    16'd37895: out <= 16'hFFCB;
    16'd37896: out <= 16'hFF19;    16'd37897: out <= 16'h00F0;    16'd37898: out <= 16'hFE31;    16'd37899: out <= 16'h036A;
    16'd37900: out <= 16'h00F6;    16'd37901: out <= 16'h02A7;    16'd37902: out <= 16'h031D;    16'd37903: out <= 16'hFAC7;
    16'd37904: out <= 16'hFC34;    16'd37905: out <= 16'h00A9;    16'd37906: out <= 16'hFEEC;    16'd37907: out <= 16'h009E;
    16'd37908: out <= 16'hFB2B;    16'd37909: out <= 16'h0254;    16'd37910: out <= 16'hFFD6;    16'd37911: out <= 16'hFA16;
    16'd37912: out <= 16'h005A;    16'd37913: out <= 16'hFFFE;    16'd37914: out <= 16'h07A7;    16'd37915: out <= 16'h01CC;
    16'd37916: out <= 16'h03D1;    16'd37917: out <= 16'hFFA3;    16'd37918: out <= 16'h0620;    16'd37919: out <= 16'h0340;
    16'd37920: out <= 16'hFDC7;    16'd37921: out <= 16'h0C93;    16'd37922: out <= 16'h09A9;    16'd37923: out <= 16'h09E3;
    16'd37924: out <= 16'hFFC4;    16'd37925: out <= 16'h048B;    16'd37926: out <= 16'h085B;    16'd37927: out <= 16'h0210;
    16'd37928: out <= 16'h01DA;    16'd37929: out <= 16'h0617;    16'd37930: out <= 16'h0675;    16'd37931: out <= 16'h02EE;
    16'd37932: out <= 16'h049B;    16'd37933: out <= 16'hFF8F;    16'd37934: out <= 16'h0076;    16'd37935: out <= 16'h019B;
    16'd37936: out <= 16'h0626;    16'd37937: out <= 16'h022D;    16'd37938: out <= 16'h092F;    16'd37939: out <= 16'h02C6;
    16'd37940: out <= 16'h0451;    16'd37941: out <= 16'h0445;    16'd37942: out <= 16'h018E;    16'd37943: out <= 16'h03C0;
    16'd37944: out <= 16'hFD26;    16'd37945: out <= 16'h0750;    16'd37946: out <= 16'h05D9;    16'd37947: out <= 16'h02E4;
    16'd37948: out <= 16'hFABD;    16'd37949: out <= 16'h02F0;    16'd37950: out <= 16'h082A;    16'd37951: out <= 16'h067A;
    16'd37952: out <= 16'h03C0;    16'd37953: out <= 16'h02D6;    16'd37954: out <= 16'h03CF;    16'd37955: out <= 16'h03C8;
    16'd37956: out <= 16'h03F5;    16'd37957: out <= 16'h06F2;    16'd37958: out <= 16'h0AD1;    16'd37959: out <= 16'h0459;
    16'd37960: out <= 16'h05D8;    16'd37961: out <= 16'h01B4;    16'd37962: out <= 16'hFE63;    16'd37963: out <= 16'h07C6;
    16'd37964: out <= 16'hFB30;    16'd37965: out <= 16'h0AF8;    16'd37966: out <= 16'h07C4;    16'd37967: out <= 16'h0728;
    16'd37968: out <= 16'hFDAD;    16'd37969: out <= 16'h0DAD;    16'd37970: out <= 16'h0B54;    16'd37971: out <= 16'hFC08;
    16'd37972: out <= 16'h008C;    16'd37973: out <= 16'h037E;    16'd37974: out <= 16'h056D;    16'd37975: out <= 16'h0589;
    16'd37976: out <= 16'h04F1;    16'd37977: out <= 16'h0C6C;    16'd37978: out <= 16'h0227;    16'd37979: out <= 16'h0A51;
    16'd37980: out <= 16'h018C;    16'd37981: out <= 16'h0498;    16'd37982: out <= 16'h0324;    16'd37983: out <= 16'h0452;
    16'd37984: out <= 16'h001A;    16'd37985: out <= 16'h023D;    16'd37986: out <= 16'h038B;    16'd37987: out <= 16'h0744;
    16'd37988: out <= 16'h01CD;    16'd37989: out <= 16'h0613;    16'd37990: out <= 16'hFFD8;    16'd37991: out <= 16'h0823;
    16'd37992: out <= 16'h06F1;    16'd37993: out <= 16'hFEDC;    16'd37994: out <= 16'h02BB;    16'd37995: out <= 16'h0B03;
    16'd37996: out <= 16'hFF29;    16'd37997: out <= 16'hFE57;    16'd37998: out <= 16'hFF46;    16'd37999: out <= 16'h02EE;
    16'd38000: out <= 16'hFC43;    16'd38001: out <= 16'h0A54;    16'd38002: out <= 16'h044C;    16'd38003: out <= 16'h0846;
    16'd38004: out <= 16'hFEE5;    16'd38005: out <= 16'hFD09;    16'd38006: out <= 16'hF3BE;    16'd38007: out <= 16'hFEF0;
    16'd38008: out <= 16'hFB12;    16'd38009: out <= 16'h0361;    16'd38010: out <= 16'h080C;    16'd38011: out <= 16'h0429;
    16'd38012: out <= 16'h0327;    16'd38013: out <= 16'hFB78;    16'd38014: out <= 16'h01A3;    16'd38015: out <= 16'h0680;
    16'd38016: out <= 16'h03AB;    16'd38017: out <= 16'hFF5C;    16'd38018: out <= 16'hFF29;    16'd38019: out <= 16'h000F;
    16'd38020: out <= 16'h030C;    16'd38021: out <= 16'hFF77;    16'd38022: out <= 16'h01DD;    16'd38023: out <= 16'hFE18;
    16'd38024: out <= 16'h062F;    16'd38025: out <= 16'hFB62;    16'd38026: out <= 16'h018E;    16'd38027: out <= 16'h04F1;
    16'd38028: out <= 16'h05A1;    16'd38029: out <= 16'h01F0;    16'd38030: out <= 16'h085A;    16'd38031: out <= 16'h04E8;
    16'd38032: out <= 16'hFD04;    16'd38033: out <= 16'h0744;    16'd38034: out <= 16'h06B1;    16'd38035: out <= 16'hFCAA;
    16'd38036: out <= 16'h0C5F;    16'd38037: out <= 16'h03CA;    16'd38038: out <= 16'h0019;    16'd38039: out <= 16'hFE33;
    16'd38040: out <= 16'h03D9;    16'd38041: out <= 16'h0799;    16'd38042: out <= 16'h0B1D;    16'd38043: out <= 16'h050E;
    16'd38044: out <= 16'h0065;    16'd38045: out <= 16'h040A;    16'd38046: out <= 16'h0698;    16'd38047: out <= 16'h03BB;
    16'd38048: out <= 16'hFD8E;    16'd38049: out <= 16'h04FD;    16'd38050: out <= 16'hFEE1;    16'd38051: out <= 16'h0A46;
    16'd38052: out <= 16'h074B;    16'd38053: out <= 16'h0120;    16'd38054: out <= 16'h02F7;    16'd38055: out <= 16'h014D;
    16'd38056: out <= 16'h0130;    16'd38057: out <= 16'h0246;    16'd38058: out <= 16'h0646;    16'd38059: out <= 16'h05DD;
    16'd38060: out <= 16'h062C;    16'd38061: out <= 16'h031A;    16'd38062: out <= 16'h02D4;    16'd38063: out <= 16'h079E;
    16'd38064: out <= 16'h079B;    16'd38065: out <= 16'hF909;    16'd38066: out <= 16'h0433;    16'd38067: out <= 16'h09F3;
    16'd38068: out <= 16'h02F0;    16'd38069: out <= 16'h0071;    16'd38070: out <= 16'h0830;    16'd38071: out <= 16'h0813;
    16'd38072: out <= 16'h0538;    16'd38073: out <= 16'h00BC;    16'd38074: out <= 16'h05B2;    16'd38075: out <= 16'h03F0;
    16'd38076: out <= 16'h02BE;    16'd38077: out <= 16'h0477;    16'd38078: out <= 16'hFE9F;    16'd38079: out <= 16'h0009;
    16'd38080: out <= 16'h00FB;    16'd38081: out <= 16'hFBC9;    16'd38082: out <= 16'hFF37;    16'd38083: out <= 16'h045E;
    16'd38084: out <= 16'hFE0F;    16'd38085: out <= 16'h0842;    16'd38086: out <= 16'h00A5;    16'd38087: out <= 16'h030C;
    16'd38088: out <= 16'h014D;    16'd38089: out <= 16'hFE40;    16'd38090: out <= 16'h032B;    16'd38091: out <= 16'h0129;
    16'd38092: out <= 16'h0A88;    16'd38093: out <= 16'h039D;    16'd38094: out <= 16'h0328;    16'd38095: out <= 16'h0346;
    16'd38096: out <= 16'h01C0;    16'd38097: out <= 16'h0490;    16'd38098: out <= 16'h0636;    16'd38099: out <= 16'h0288;
    16'd38100: out <= 16'h04F8;    16'd38101: out <= 16'hFD58;    16'd38102: out <= 16'hFE37;    16'd38103: out <= 16'hFF3B;
    16'd38104: out <= 16'h0014;    16'd38105: out <= 16'h032A;    16'd38106: out <= 16'h07B1;    16'd38107: out <= 16'h0648;
    16'd38108: out <= 16'h0089;    16'd38109: out <= 16'h0781;    16'd38110: out <= 16'h078C;    16'd38111: out <= 16'h006B;
    16'd38112: out <= 16'h056E;    16'd38113: out <= 16'h0126;    16'd38114: out <= 16'h0173;    16'd38115: out <= 16'hFE67;
    16'd38116: out <= 16'h04B8;    16'd38117: out <= 16'hFF6B;    16'd38118: out <= 16'h00DE;    16'd38119: out <= 16'hFF34;
    16'd38120: out <= 16'h0327;    16'd38121: out <= 16'h04F9;    16'd38122: out <= 16'h02AB;    16'd38123: out <= 16'hFB36;
    16'd38124: out <= 16'h0935;    16'd38125: out <= 16'h03FA;    16'd38126: out <= 16'h01A1;    16'd38127: out <= 16'hFF1B;
    16'd38128: out <= 16'h02EB;    16'd38129: out <= 16'hFE71;    16'd38130: out <= 16'hFBCE;    16'd38131: out <= 16'h04B4;
    16'd38132: out <= 16'hFD25;    16'd38133: out <= 16'h01DA;    16'd38134: out <= 16'hF792;    16'd38135: out <= 16'hFCB8;
    16'd38136: out <= 16'h0200;    16'd38137: out <= 16'h02B1;    16'd38138: out <= 16'h0418;    16'd38139: out <= 16'h0499;
    16'd38140: out <= 16'h0518;    16'd38141: out <= 16'hFAD3;    16'd38142: out <= 16'h0360;    16'd38143: out <= 16'hFF33;
    16'd38144: out <= 16'h0924;    16'd38145: out <= 16'hFBD8;    16'd38146: out <= 16'hF82B;    16'd38147: out <= 16'h068D;
    16'd38148: out <= 16'h01D9;    16'd38149: out <= 16'hFE11;    16'd38150: out <= 16'h05BB;    16'd38151: out <= 16'hFF0A;
    16'd38152: out <= 16'hFF3B;    16'd38153: out <= 16'hFEC2;    16'd38154: out <= 16'hF85B;    16'd38155: out <= 16'hFE1A;
    16'd38156: out <= 16'h034C;    16'd38157: out <= 16'h04B3;    16'd38158: out <= 16'hFAA7;    16'd38159: out <= 16'hFFD6;
    16'd38160: out <= 16'hF932;    16'd38161: out <= 16'h058C;    16'd38162: out <= 16'h038B;    16'd38163: out <= 16'h00BC;
    16'd38164: out <= 16'hFF7F;    16'd38165: out <= 16'hFC4E;    16'd38166: out <= 16'hFD95;    16'd38167: out <= 16'hF378;
    16'd38168: out <= 16'hFC45;    16'd38169: out <= 16'hFE81;    16'd38170: out <= 16'h00E5;    16'd38171: out <= 16'h0272;
    16'd38172: out <= 16'h0520;    16'd38173: out <= 16'h0605;    16'd38174: out <= 16'h04A1;    16'd38175: out <= 16'h039E;
    16'd38176: out <= 16'hFE17;    16'd38177: out <= 16'h03E4;    16'd38178: out <= 16'h02F9;    16'd38179: out <= 16'h074C;
    16'd38180: out <= 16'h031B;    16'd38181: out <= 16'h033B;    16'd38182: out <= 16'h0022;    16'd38183: out <= 16'h0063;
    16'd38184: out <= 16'h05CD;    16'd38185: out <= 16'h0074;    16'd38186: out <= 16'h009E;    16'd38187: out <= 16'hFE48;
    16'd38188: out <= 16'h0A49;    16'd38189: out <= 16'h0797;    16'd38190: out <= 16'h0040;    16'd38191: out <= 16'h02E5;
    16'd38192: out <= 16'h0875;    16'd38193: out <= 16'h05DF;    16'd38194: out <= 16'h0547;    16'd38195: out <= 16'h041C;
    16'd38196: out <= 16'h03F8;    16'd38197: out <= 16'h00B7;    16'd38198: out <= 16'h0504;    16'd38199: out <= 16'h04C9;
    16'd38200: out <= 16'h075D;    16'd38201: out <= 16'h0C62;    16'd38202: out <= 16'h025A;    16'd38203: out <= 16'h0623;
    16'd38204: out <= 16'hFFB9;    16'd38205: out <= 16'h08FD;    16'd38206: out <= 16'h0190;    16'd38207: out <= 16'h0222;
    16'd38208: out <= 16'h05B5;    16'd38209: out <= 16'h00FA;    16'd38210: out <= 16'h0087;    16'd38211: out <= 16'h0105;
    16'd38212: out <= 16'h0136;    16'd38213: out <= 16'h04C0;    16'd38214: out <= 16'h0988;    16'd38215: out <= 16'h08A4;
    16'd38216: out <= 16'h005C;    16'd38217: out <= 16'h0B1B;    16'd38218: out <= 16'hFEE3;    16'd38219: out <= 16'hFDCF;
    16'd38220: out <= 16'h0652;    16'd38221: out <= 16'h057E;    16'd38222: out <= 16'h0270;    16'd38223: out <= 16'h0250;
    16'd38224: out <= 16'h04FF;    16'd38225: out <= 16'h07AF;    16'd38226: out <= 16'h02E0;    16'd38227: out <= 16'h0337;
    16'd38228: out <= 16'h06E9;    16'd38229: out <= 16'h010C;    16'd38230: out <= 16'h0500;    16'd38231: out <= 16'hFDC3;
    16'd38232: out <= 16'h0703;    16'd38233: out <= 16'hFEFF;    16'd38234: out <= 16'h01A4;    16'd38235: out <= 16'h0577;
    16'd38236: out <= 16'h059F;    16'd38237: out <= 16'h0137;    16'd38238: out <= 16'h039B;    16'd38239: out <= 16'h0914;
    16'd38240: out <= 16'h047E;    16'd38241: out <= 16'h01A4;    16'd38242: out <= 16'h066A;    16'd38243: out <= 16'h01C2;
    16'd38244: out <= 16'h0820;    16'd38245: out <= 16'h02DB;    16'd38246: out <= 16'h05EE;    16'd38247: out <= 16'h032A;
    16'd38248: out <= 16'hFFF8;    16'd38249: out <= 16'h06FD;    16'd38250: out <= 16'h0DE9;    16'd38251: out <= 16'h0081;
    16'd38252: out <= 16'h0802;    16'd38253: out <= 16'h0385;    16'd38254: out <= 16'hFD2F;    16'd38255: out <= 16'h03C9;
    16'd38256: out <= 16'h0094;    16'd38257: out <= 16'hFBEA;    16'd38258: out <= 16'h00BB;    16'd38259: out <= 16'h0668;
    16'd38260: out <= 16'h0035;    16'd38261: out <= 16'h026B;    16'd38262: out <= 16'hFBC3;    16'd38263: out <= 16'hF844;
    16'd38264: out <= 16'h0188;    16'd38265: out <= 16'hFF5F;    16'd38266: out <= 16'hFB35;    16'd38267: out <= 16'h05E5;
    16'd38268: out <= 16'h042E;    16'd38269: out <= 16'h0207;    16'd38270: out <= 16'h051C;    16'd38271: out <= 16'h02AA;
    16'd38272: out <= 16'h047D;    16'd38273: out <= 16'hFF8A;    16'd38274: out <= 16'h03B4;    16'd38275: out <= 16'h03B5;
    16'd38276: out <= 16'hF9CA;    16'd38277: out <= 16'h04F8;    16'd38278: out <= 16'h04F0;    16'd38279: out <= 16'h032F;
    16'd38280: out <= 16'h02A5;    16'd38281: out <= 16'h0463;    16'd38282: out <= 16'hFEC5;    16'd38283: out <= 16'h0A55;
    16'd38284: out <= 16'h0875;    16'd38285: out <= 16'h0939;    16'd38286: out <= 16'h01A1;    16'd38287: out <= 16'h0442;
    16'd38288: out <= 16'h08CE;    16'd38289: out <= 16'h09C8;    16'd38290: out <= 16'hFFE5;    16'd38291: out <= 16'h0162;
    16'd38292: out <= 16'h055D;    16'd38293: out <= 16'h0087;    16'd38294: out <= 16'h022B;    16'd38295: out <= 16'hFCF7;
    16'd38296: out <= 16'h0106;    16'd38297: out <= 16'h0475;    16'd38298: out <= 16'h0A3E;    16'd38299: out <= 16'h03A2;
    16'd38300: out <= 16'h066D;    16'd38301: out <= 16'hFFB9;    16'd38302: out <= 16'hFEE4;    16'd38303: out <= 16'h05F1;
    16'd38304: out <= 16'h08F8;    16'd38305: out <= 16'h04CC;    16'd38306: out <= 16'hFEFA;    16'd38307: out <= 16'h01F7;
    16'd38308: out <= 16'hFFDD;    16'd38309: out <= 16'h0020;    16'd38310: out <= 16'h0784;    16'd38311: out <= 16'h0455;
    16'd38312: out <= 16'h00BF;    16'd38313: out <= 16'h0721;    16'd38314: out <= 16'h01D9;    16'd38315: out <= 16'h03D8;
    16'd38316: out <= 16'h0169;    16'd38317: out <= 16'h0455;    16'd38318: out <= 16'h0A95;    16'd38319: out <= 16'h0235;
    16'd38320: out <= 16'h0ACD;    16'd38321: out <= 16'h0710;    16'd38322: out <= 16'h086F;    16'd38323: out <= 16'h0264;
    16'd38324: out <= 16'h04DF;    16'd38325: out <= 16'h057A;    16'd38326: out <= 16'h0235;    16'd38327: out <= 16'h0154;
    16'd38328: out <= 16'h0E1C;    16'd38329: out <= 16'h0A38;    16'd38330: out <= 16'h02A3;    16'd38331: out <= 16'h0496;
    16'd38332: out <= 16'hFFCB;    16'd38333: out <= 16'h01CF;    16'd38334: out <= 16'h01DA;    16'd38335: out <= 16'h03DB;
    16'd38336: out <= 16'h03B2;    16'd38337: out <= 16'h0077;    16'd38338: out <= 16'h0044;    16'd38339: out <= 16'h03B6;
    16'd38340: out <= 16'hFF6F;    16'd38341: out <= 16'hFF6C;    16'd38342: out <= 16'h05C9;    16'd38343: out <= 16'h04B2;
    16'd38344: out <= 16'hFCFA;    16'd38345: out <= 16'h0179;    16'd38346: out <= 16'h000D;    16'd38347: out <= 16'h0011;
    16'd38348: out <= 16'h0502;    16'd38349: out <= 16'h0178;    16'd38350: out <= 16'h070A;    16'd38351: out <= 16'h0585;
    16'd38352: out <= 16'h0220;    16'd38353: out <= 16'h02A2;    16'd38354: out <= 16'hFFF5;    16'd38355: out <= 16'h05EE;
    16'd38356: out <= 16'h082E;    16'd38357: out <= 16'h056E;    16'd38358: out <= 16'h01B0;    16'd38359: out <= 16'hFDDB;
    16'd38360: out <= 16'h0840;    16'd38361: out <= 16'h01F5;    16'd38362: out <= 16'hFAE9;    16'd38363: out <= 16'h071E;
    16'd38364: out <= 16'h07CA;    16'd38365: out <= 16'h0786;    16'd38366: out <= 16'h046A;    16'd38367: out <= 16'h0403;
    16'd38368: out <= 16'h07C3;    16'd38369: out <= 16'h007F;    16'd38370: out <= 16'h0A02;    16'd38371: out <= 16'h01FD;
    16'd38372: out <= 16'h060F;    16'd38373: out <= 16'h03FF;    16'd38374: out <= 16'h063C;    16'd38375: out <= 16'hFA8B;
    16'd38376: out <= 16'hFCA4;    16'd38377: out <= 16'h0017;    16'd38378: out <= 16'h00EC;    16'd38379: out <= 16'hFDDF;
    16'd38380: out <= 16'h04B7;    16'd38381: out <= 16'h0749;    16'd38382: out <= 16'hFDA2;    16'd38383: out <= 16'h02F8;
    16'd38384: out <= 16'hFA80;    16'd38385: out <= 16'hFFA2;    16'd38386: out <= 16'h00A4;    16'd38387: out <= 16'hFC02;
    16'd38388: out <= 16'h0117;    16'd38389: out <= 16'h0385;    16'd38390: out <= 16'hFA63;    16'd38391: out <= 16'h004E;
    16'd38392: out <= 16'hFBE8;    16'd38393: out <= 16'hF9E8;    16'd38394: out <= 16'hFFCC;    16'd38395: out <= 16'hFB7D;
    16'd38396: out <= 16'hFC51;    16'd38397: out <= 16'h0372;    16'd38398: out <= 16'hFF67;    16'd38399: out <= 16'hFB05;
    16'd38400: out <= 16'hFDCE;    16'd38401: out <= 16'h012C;    16'd38402: out <= 16'hFFB8;    16'd38403: out <= 16'hFA7F;
    16'd38404: out <= 16'h0325;    16'd38405: out <= 16'hFC0E;    16'd38406: out <= 16'h036B;    16'd38407: out <= 16'h0025;
    16'd38408: out <= 16'hF7B4;    16'd38409: out <= 16'hFF91;    16'd38410: out <= 16'h0082;    16'd38411: out <= 16'hFE73;
    16'd38412: out <= 16'hF734;    16'd38413: out <= 16'h006C;    16'd38414: out <= 16'hFCA0;    16'd38415: out <= 16'hFE8D;
    16'd38416: out <= 16'hFF88;    16'd38417: out <= 16'hF852;    16'd38418: out <= 16'h0690;    16'd38419: out <= 16'hF956;
    16'd38420: out <= 16'h021F;    16'd38421: out <= 16'hFF1C;    16'd38422: out <= 16'hFF63;    16'd38423: out <= 16'h00AE;
    16'd38424: out <= 16'hFA61;    16'd38425: out <= 16'hFD41;    16'd38426: out <= 16'h0605;    16'd38427: out <= 16'h02D0;
    16'd38428: out <= 16'h02F4;    16'd38429: out <= 16'h062E;    16'd38430: out <= 16'hFC65;    16'd38431: out <= 16'h071D;
    16'd38432: out <= 16'hFFA3;    16'd38433: out <= 16'h020E;    16'd38434: out <= 16'h0475;    16'd38435: out <= 16'h05BB;
    16'd38436: out <= 16'h070F;    16'd38437: out <= 16'h091C;    16'd38438: out <= 16'hFD90;    16'd38439: out <= 16'h0623;
    16'd38440: out <= 16'hFFE9;    16'd38441: out <= 16'h04DA;    16'd38442: out <= 16'h0C88;    16'd38443: out <= 16'h00DD;
    16'd38444: out <= 16'h03FD;    16'd38445: out <= 16'h000A;    16'd38446: out <= 16'h09E0;    16'd38447: out <= 16'h0602;
    16'd38448: out <= 16'h0C2F;    16'd38449: out <= 16'h0C45;    16'd38450: out <= 16'h085A;    16'd38451: out <= 16'h025B;
    16'd38452: out <= 16'h05DA;    16'd38453: out <= 16'hFE75;    16'd38454: out <= 16'h07BE;    16'd38455: out <= 16'h0362;
    16'd38456: out <= 16'hFF55;    16'd38457: out <= 16'h06CC;    16'd38458: out <= 16'h0090;    16'd38459: out <= 16'hFDF3;
    16'd38460: out <= 16'h0524;    16'd38461: out <= 16'h0668;    16'd38462: out <= 16'h0539;    16'd38463: out <= 16'h0CA9;
    16'd38464: out <= 16'h02A8;    16'd38465: out <= 16'h0774;    16'd38466: out <= 16'h02B8;    16'd38467: out <= 16'h05B1;
    16'd38468: out <= 16'h063D;    16'd38469: out <= 16'h0594;    16'd38470: out <= 16'h0239;    16'd38471: out <= 16'h07B1;
    16'd38472: out <= 16'h03E3;    16'd38473: out <= 16'hFF34;    16'd38474: out <= 16'hFE9C;    16'd38475: out <= 16'h06D2;
    16'd38476: out <= 16'h02A9;    16'd38477: out <= 16'hF9BE;    16'd38478: out <= 16'h0121;    16'd38479: out <= 16'hFB8C;
    16'd38480: out <= 16'h01EB;    16'd38481: out <= 16'h06B8;    16'd38482: out <= 16'h00A1;    16'd38483: out <= 16'hF984;
    16'd38484: out <= 16'h043A;    16'd38485: out <= 16'h0647;    16'd38486: out <= 16'h073A;    16'd38487: out <= 16'h043A;
    16'd38488: out <= 16'h042E;    16'd38489: out <= 16'h09F1;    16'd38490: out <= 16'h02F8;    16'd38491: out <= 16'h00F4;
    16'd38492: out <= 16'h064B;    16'd38493: out <= 16'h03FA;    16'd38494: out <= 16'h0458;    16'd38495: out <= 16'h05E2;
    16'd38496: out <= 16'h020E;    16'd38497: out <= 16'h00A7;    16'd38498: out <= 16'h07AD;    16'd38499: out <= 16'h0809;
    16'd38500: out <= 16'h0667;    16'd38501: out <= 16'h01AF;    16'd38502: out <= 16'h03AD;    16'd38503: out <= 16'h05DD;
    16'd38504: out <= 16'h0482;    16'd38505: out <= 16'h04FE;    16'd38506: out <= 16'h0678;    16'd38507: out <= 16'h02B8;
    16'd38508: out <= 16'hFED1;    16'd38509: out <= 16'h049E;    16'd38510: out <= 16'h012B;    16'd38511: out <= 16'hFF35;
    16'd38512: out <= 16'hFB1B;    16'd38513: out <= 16'h048E;    16'd38514: out <= 16'h0267;    16'd38515: out <= 16'h004C;
    16'd38516: out <= 16'hFD67;    16'd38517: out <= 16'h0053;    16'd38518: out <= 16'h07A1;    16'd38519: out <= 16'hFFBD;
    16'd38520: out <= 16'h058B;    16'd38521: out <= 16'h039F;    16'd38522: out <= 16'hFED3;    16'd38523: out <= 16'h0521;
    16'd38524: out <= 16'h01E3;    16'd38525: out <= 16'h0699;    16'd38526: out <= 16'h079A;    16'd38527: out <= 16'h04F3;
    16'd38528: out <= 16'h0342;    16'd38529: out <= 16'hFF02;    16'd38530: out <= 16'h0985;    16'd38531: out <= 16'h050C;
    16'd38532: out <= 16'h006D;    16'd38533: out <= 16'hFFE5;    16'd38534: out <= 16'h0166;    16'd38535: out <= 16'h06EB;
    16'd38536: out <= 16'h0393;    16'd38537: out <= 16'h04DB;    16'd38538: out <= 16'h0268;    16'd38539: out <= 16'h0516;
    16'd38540: out <= 16'h0264;    16'd38541: out <= 16'h06BC;    16'd38542: out <= 16'h06ED;    16'd38543: out <= 16'h0483;
    16'd38544: out <= 16'h0645;    16'd38545: out <= 16'h031E;    16'd38546: out <= 16'h0AB5;    16'd38547: out <= 16'h046A;
    16'd38548: out <= 16'h04DC;    16'd38549: out <= 16'h0240;    16'd38550: out <= 16'h0785;    16'd38551: out <= 16'h09FC;
    16'd38552: out <= 16'h07A7;    16'd38553: out <= 16'h0C9B;    16'd38554: out <= 16'h08D0;    16'd38555: out <= 16'h0107;
    16'd38556: out <= 16'h0672;    16'd38557: out <= 16'h05A6;    16'd38558: out <= 16'h00DF;    16'd38559: out <= 16'h03F2;
    16'd38560: out <= 16'hFF79;    16'd38561: out <= 16'hFEDD;    16'd38562: out <= 16'h0AD7;    16'd38563: out <= 16'hFEC0;
    16'd38564: out <= 16'h04C7;    16'd38565: out <= 16'h02B5;    16'd38566: out <= 16'hFD60;    16'd38567: out <= 16'h0134;
    16'd38568: out <= 16'h08E7;    16'd38569: out <= 16'hFF57;    16'd38570: out <= 16'h02F5;    16'd38571: out <= 16'hFCF6;
    16'd38572: out <= 16'hFD04;    16'd38573: out <= 16'h04D1;    16'd38574: out <= 16'h01E7;    16'd38575: out <= 16'h044D;
    16'd38576: out <= 16'h046E;    16'd38577: out <= 16'h09AF;    16'd38578: out <= 16'h091C;    16'd38579: out <= 16'h04B6;
    16'd38580: out <= 16'h0379;    16'd38581: out <= 16'h0A5F;    16'd38582: out <= 16'h02E2;    16'd38583: out <= 16'h0753;
    16'd38584: out <= 16'h0569;    16'd38585: out <= 16'h03A6;    16'd38586: out <= 16'h051C;    16'd38587: out <= 16'hFFF5;
    16'd38588: out <= 16'hFD12;    16'd38589: out <= 16'h02E6;    16'd38590: out <= 16'h0412;    16'd38591: out <= 16'h063E;
    16'd38592: out <= 16'h01B5;    16'd38593: out <= 16'h05B1;    16'd38594: out <= 16'hFF95;    16'd38595: out <= 16'h02DF;
    16'd38596: out <= 16'h0C77;    16'd38597: out <= 16'h06F6;    16'd38598: out <= 16'h01F7;    16'd38599: out <= 16'h03E5;
    16'd38600: out <= 16'h0105;    16'd38601: out <= 16'hFEA5;    16'd38602: out <= 16'h0966;    16'd38603: out <= 16'h01AD;
    16'd38604: out <= 16'h0037;    16'd38605: out <= 16'h05C2;    16'd38606: out <= 16'h0594;    16'd38607: out <= 16'h034C;
    16'd38608: out <= 16'h08D3;    16'd38609: out <= 16'h0876;    16'd38610: out <= 16'hFF43;    16'd38611: out <= 16'h0C86;
    16'd38612: out <= 16'h01CC;    16'd38613: out <= 16'hFF17;    16'd38614: out <= 16'hF77B;    16'd38615: out <= 16'h033B;
    16'd38616: out <= 16'h04EE;    16'd38617: out <= 16'h03C9;    16'd38618: out <= 16'h027A;    16'd38619: out <= 16'h019C;
    16'd38620: out <= 16'h01B1;    16'd38621: out <= 16'h0A0B;    16'd38622: out <= 16'h05EA;    16'd38623: out <= 16'h03D4;
    16'd38624: out <= 16'h04E7;    16'd38625: out <= 16'h029E;    16'd38626: out <= 16'h007C;    16'd38627: out <= 16'h032E;
    16'd38628: out <= 16'h0735;    16'd38629: out <= 16'hFF61;    16'd38630: out <= 16'h02CC;    16'd38631: out <= 16'hFD82;
    16'd38632: out <= 16'hFDBF;    16'd38633: out <= 16'hF8FC;    16'd38634: out <= 16'h0636;    16'd38635: out <= 16'h003C;
    16'd38636: out <= 16'hFC56;    16'd38637: out <= 16'hF9DA;    16'd38638: out <= 16'hF88B;    16'd38639: out <= 16'hFBE4;
    16'd38640: out <= 16'hF914;    16'd38641: out <= 16'hFBDF;    16'd38642: out <= 16'h00B8;    16'd38643: out <= 16'hFEC4;
    16'd38644: out <= 16'hFBF4;    16'd38645: out <= 16'h0193;    16'd38646: out <= 16'hFAC8;    16'd38647: out <= 16'h028A;
    16'd38648: out <= 16'h03BB;    16'd38649: out <= 16'h0295;    16'd38650: out <= 16'hFFCD;    16'd38651: out <= 16'h03C4;
    16'd38652: out <= 16'h0115;    16'd38653: out <= 16'hFC49;    16'd38654: out <= 16'hFE6B;    16'd38655: out <= 16'h03A6;
    16'd38656: out <= 16'h02B4;    16'd38657: out <= 16'hFC2D;    16'd38658: out <= 16'hFD51;    16'd38659: out <= 16'hFED3;
    16'd38660: out <= 16'h021C;    16'd38661: out <= 16'hFB11;    16'd38662: out <= 16'hFC01;    16'd38663: out <= 16'h03B2;
    16'd38664: out <= 16'hFC1D;    16'd38665: out <= 16'h04D1;    16'd38666: out <= 16'h0038;    16'd38667: out <= 16'hF5BB;
    16'd38668: out <= 16'h0200;    16'd38669: out <= 16'hFAC2;    16'd38670: out <= 16'hFE78;    16'd38671: out <= 16'hFB2B;
    16'd38672: out <= 16'hFC45;    16'd38673: out <= 16'hFB91;    16'd38674: out <= 16'hFF8C;    16'd38675: out <= 16'h021F;
    16'd38676: out <= 16'hFA93;    16'd38677: out <= 16'hFA02;    16'd38678: out <= 16'h01ED;    16'd38679: out <= 16'h044F;
    16'd38680: out <= 16'h014D;    16'd38681: out <= 16'h0692;    16'd38682: out <= 16'hFC3A;    16'd38683: out <= 16'h0690;
    16'd38684: out <= 16'h0397;    16'd38685: out <= 16'h03F3;    16'd38686: out <= 16'h04A5;    16'd38687: out <= 16'h04E8;
    16'd38688: out <= 16'hFD65;    16'd38689: out <= 16'h040D;    16'd38690: out <= 16'h053F;    16'd38691: out <= 16'h0026;
    16'd38692: out <= 16'h00D5;    16'd38693: out <= 16'h0957;    16'd38694: out <= 16'h0163;    16'd38695: out <= 16'h0071;
    16'd38696: out <= 16'h04A2;    16'd38697: out <= 16'h026F;    16'd38698: out <= 16'h0245;    16'd38699: out <= 16'h00AB;
    16'd38700: out <= 16'h0599;    16'd38701: out <= 16'hFB3C;    16'd38702: out <= 16'h048A;    16'd38703: out <= 16'h05A4;
    16'd38704: out <= 16'h0746;    16'd38705: out <= 16'h059D;    16'd38706: out <= 16'h08F5;    16'd38707: out <= 16'hFE5E;
    16'd38708: out <= 16'h038B;    16'd38709: out <= 16'h004A;    16'd38710: out <= 16'h03B3;    16'd38711: out <= 16'hFE7A;
    16'd38712: out <= 16'hFBDD;    16'd38713: out <= 16'h0949;    16'd38714: out <= 16'h098A;    16'd38715: out <= 16'hFFC8;
    16'd38716: out <= 16'h042A;    16'd38717: out <= 16'h0110;    16'd38718: out <= 16'hFFF6;    16'd38719: out <= 16'hFE74;
    16'd38720: out <= 16'h037B;    16'd38721: out <= 16'h0577;    16'd38722: out <= 16'h0A0A;    16'd38723: out <= 16'h05B6;
    16'd38724: out <= 16'h077C;    16'd38725: out <= 16'h0842;    16'd38726: out <= 16'h0195;    16'd38727: out <= 16'h06DF;
    16'd38728: out <= 16'h02AC;    16'd38729: out <= 16'h0889;    16'd38730: out <= 16'h039E;    16'd38731: out <= 16'hFB39;
    16'd38732: out <= 16'hFF61;    16'd38733: out <= 16'h055F;    16'd38734: out <= 16'h0102;    16'd38735: out <= 16'hFFC6;
    16'd38736: out <= 16'h0CEA;    16'd38737: out <= 16'h0446;    16'd38738: out <= 16'hFF9C;    16'd38739: out <= 16'h0507;
    16'd38740: out <= 16'h05A9;    16'd38741: out <= 16'h03D8;    16'd38742: out <= 16'h0A70;    16'd38743: out <= 16'h0404;
    16'd38744: out <= 16'hFFB4;    16'd38745: out <= 16'h05F9;    16'd38746: out <= 16'h0787;    16'd38747: out <= 16'h01AC;
    16'd38748: out <= 16'h0ABD;    16'd38749: out <= 16'h0105;    16'd38750: out <= 16'h0736;    16'd38751: out <= 16'h03FD;
    16'd38752: out <= 16'h0780;    16'd38753: out <= 16'h0747;    16'd38754: out <= 16'h0AEB;    16'd38755: out <= 16'h021E;
    16'd38756: out <= 16'h0303;    16'd38757: out <= 16'h0596;    16'd38758: out <= 16'h0A66;    16'd38759: out <= 16'h0929;
    16'd38760: out <= 16'h0323;    16'd38761: out <= 16'hFD2B;    16'd38762: out <= 16'hFE01;    16'd38763: out <= 16'hFFDA;
    16'd38764: out <= 16'h05ED;    16'd38765: out <= 16'h01E1;    16'd38766: out <= 16'hF9B3;    16'd38767: out <= 16'h024D;
    16'd38768: out <= 16'h0373;    16'd38769: out <= 16'h055A;    16'd38770: out <= 16'h03ED;    16'd38771: out <= 16'h008D;
    16'd38772: out <= 16'hFA62;    16'd38773: out <= 16'hF9F8;    16'd38774: out <= 16'hFF24;    16'd38775: out <= 16'h058F;
    16'd38776: out <= 16'h00AB;    16'd38777: out <= 16'hFBAF;    16'd38778: out <= 16'h0300;    16'd38779: out <= 16'h0739;
    16'd38780: out <= 16'h0873;    16'd38781: out <= 16'hFF73;    16'd38782: out <= 16'h00D6;    16'd38783: out <= 16'h0355;
    16'd38784: out <= 16'hFFC0;    16'd38785: out <= 16'h05A0;    16'd38786: out <= 16'h0710;    16'd38787: out <= 16'h0256;
    16'd38788: out <= 16'h0994;    16'd38789: out <= 16'h05C6;    16'd38790: out <= 16'h0758;    16'd38791: out <= 16'h06C9;
    16'd38792: out <= 16'h0BF5;    16'd38793: out <= 16'h08C2;    16'd38794: out <= 16'h0515;    16'd38795: out <= 16'h07A2;
    16'd38796: out <= 16'h0252;    16'd38797: out <= 16'h0318;    16'd38798: out <= 16'h087F;    16'd38799: out <= 16'h064D;
    16'd38800: out <= 16'h0075;    16'd38801: out <= 16'h0576;    16'd38802: out <= 16'h0029;    16'd38803: out <= 16'h0A38;
    16'd38804: out <= 16'h08BC;    16'd38805: out <= 16'h0897;    16'd38806: out <= 16'h02BC;    16'd38807: out <= 16'h02EB;
    16'd38808: out <= 16'hFED2;    16'd38809: out <= 16'h011A;    16'd38810: out <= 16'hFD40;    16'd38811: out <= 16'h096B;
    16'd38812: out <= 16'h02BB;    16'd38813: out <= 16'h00D1;    16'd38814: out <= 16'h099A;    16'd38815: out <= 16'h0958;
    16'd38816: out <= 16'h0189;    16'd38817: out <= 16'h026E;    16'd38818: out <= 16'h062F;    16'd38819: out <= 16'h09AF;
    16'd38820: out <= 16'h08B1;    16'd38821: out <= 16'h08FD;    16'd38822: out <= 16'h05C3;    16'd38823: out <= 16'h060B;
    16'd38824: out <= 16'hFC88;    16'd38825: out <= 16'h00C0;    16'd38826: out <= 16'hFBF9;    16'd38827: out <= 16'h0B58;
    16'd38828: out <= 16'hFB77;    16'd38829: out <= 16'h01A2;    16'd38830: out <= 16'hFDD0;    16'd38831: out <= 16'h0705;
    16'd38832: out <= 16'h06A3;    16'd38833: out <= 16'h01D7;    16'd38834: out <= 16'h0517;    16'd38835: out <= 16'hFF1E;
    16'd38836: out <= 16'h0597;    16'd38837: out <= 16'h03F2;    16'd38838: out <= 16'h07A4;    16'd38839: out <= 16'h04C8;
    16'd38840: out <= 16'h04DD;    16'd38841: out <= 16'h00B4;    16'd38842: out <= 16'hFD43;    16'd38843: out <= 16'h06CF;
    16'd38844: out <= 16'h0180;    16'd38845: out <= 16'h0340;    16'd38846: out <= 16'h03E3;    16'd38847: out <= 16'h00F2;
    16'd38848: out <= 16'hFE34;    16'd38849: out <= 16'hFC16;    16'd38850: out <= 16'h071C;    16'd38851: out <= 16'h075F;
    16'd38852: out <= 16'h0749;    16'd38853: out <= 16'h04B3;    16'd38854: out <= 16'hFFDE;    16'd38855: out <= 16'h05ED;
    16'd38856: out <= 16'h094C;    16'd38857: out <= 16'h0703;    16'd38858: out <= 16'h02B6;    16'd38859: out <= 16'h0352;
    16'd38860: out <= 16'h0476;    16'd38861: out <= 16'hFB13;    16'd38862: out <= 16'h0081;    16'd38863: out <= 16'h0545;
    16'd38864: out <= 16'h0270;    16'd38865: out <= 16'h018D;    16'd38866: out <= 16'h00E8;    16'd38867: out <= 16'h0495;
    16'd38868: out <= 16'hFDDA;    16'd38869: out <= 16'hFE37;    16'd38870: out <= 16'hFE79;    16'd38871: out <= 16'h07FC;
    16'd38872: out <= 16'h0A60;    16'd38873: out <= 16'h017D;    16'd38874: out <= 16'hFCB2;    16'd38875: out <= 16'hFFBE;
    16'd38876: out <= 16'h01F5;    16'd38877: out <= 16'h0092;    16'd38878: out <= 16'h0858;    16'd38879: out <= 16'hFD6B;
    16'd38880: out <= 16'h0A63;    16'd38881: out <= 16'h00A8;    16'd38882: out <= 16'hFE0E;    16'd38883: out <= 16'h046C;
    16'd38884: out <= 16'h00DF;    16'd38885: out <= 16'h0043;    16'd38886: out <= 16'h0097;    16'd38887: out <= 16'hFECD;
    16'd38888: out <= 16'h0176;    16'd38889: out <= 16'hFBD8;    16'd38890: out <= 16'hFEC9;    16'd38891: out <= 16'h025A;
    16'd38892: out <= 16'h012F;    16'd38893: out <= 16'h042E;    16'd38894: out <= 16'hFC7D;    16'd38895: out <= 16'hFD94;
    16'd38896: out <= 16'hFBFD;    16'd38897: out <= 16'hFF26;    16'd38898: out <= 16'hFDDA;    16'd38899: out <= 16'hF820;
    16'd38900: out <= 16'h0582;    16'd38901: out <= 16'hFFC6;    16'd38902: out <= 16'h022B;    16'd38903: out <= 16'h0085;
    16'd38904: out <= 16'h0312;    16'd38905: out <= 16'h05D0;    16'd38906: out <= 16'h0431;    16'd38907: out <= 16'hFDF4;
    16'd38908: out <= 16'h00C7;    16'd38909: out <= 16'h0278;    16'd38910: out <= 16'hF846;    16'd38911: out <= 16'h00C0;
    16'd38912: out <= 16'hFCEF;    16'd38913: out <= 16'h049E;    16'd38914: out <= 16'h06A4;    16'd38915: out <= 16'h014B;
    16'd38916: out <= 16'hFDB4;    16'd38917: out <= 16'hF9EA;    16'd38918: out <= 16'hFC21;    16'd38919: out <= 16'hF9C1;
    16'd38920: out <= 16'hFE6F;    16'd38921: out <= 16'h02B2;    16'd38922: out <= 16'hFF7E;    16'd38923: out <= 16'hFF42;
    16'd38924: out <= 16'h05C8;    16'd38925: out <= 16'hFFDD;    16'd38926: out <= 16'h00CC;    16'd38927: out <= 16'hFD9B;
    16'd38928: out <= 16'hFCF7;    16'd38929: out <= 16'hFE9A;    16'd38930: out <= 16'hFDC3;    16'd38931: out <= 16'hFE6F;
    16'd38932: out <= 16'h0695;    16'd38933: out <= 16'hFC12;    16'd38934: out <= 16'h0075;    16'd38935: out <= 16'h0800;
    16'd38936: out <= 16'hF8B0;    16'd38937: out <= 16'h0112;    16'd38938: out <= 16'hFCA6;    16'd38939: out <= 16'h071A;
    16'd38940: out <= 16'h063A;    16'd38941: out <= 16'h065E;    16'd38942: out <= 16'h0368;    16'd38943: out <= 16'hFF5F;
    16'd38944: out <= 16'h0266;    16'd38945: out <= 16'h063D;    16'd38946: out <= 16'h017F;    16'd38947: out <= 16'h022B;
    16'd38948: out <= 16'h0065;    16'd38949: out <= 16'h0976;    16'd38950: out <= 16'h0A70;    16'd38951: out <= 16'h0350;
    16'd38952: out <= 16'h08AA;    16'd38953: out <= 16'h0225;    16'd38954: out <= 16'h0239;    16'd38955: out <= 16'h00E5;
    16'd38956: out <= 16'h0789;    16'd38957: out <= 16'h0476;    16'd38958: out <= 16'h019A;    16'd38959: out <= 16'h016C;
    16'd38960: out <= 16'h0124;    16'd38961: out <= 16'hFED3;    16'd38962: out <= 16'h0004;    16'd38963: out <= 16'h0287;
    16'd38964: out <= 16'hFDDE;    16'd38965: out <= 16'h0517;    16'd38966: out <= 16'h008E;    16'd38967: out <= 16'h04CB;
    16'd38968: out <= 16'h0B32;    16'd38969: out <= 16'hFC14;    16'd38970: out <= 16'h01A1;    16'd38971: out <= 16'hFDA3;
    16'd38972: out <= 16'h0A16;    16'd38973: out <= 16'h0147;    16'd38974: out <= 16'h02E8;    16'd38975: out <= 16'hFFF4;
    16'd38976: out <= 16'h05C3;    16'd38977: out <= 16'h058F;    16'd38978: out <= 16'h0725;    16'd38979: out <= 16'h0602;
    16'd38980: out <= 16'h0ACE;    16'd38981: out <= 16'hFF17;    16'd38982: out <= 16'h02C5;    16'd38983: out <= 16'h00C2;
    16'd38984: out <= 16'h0758;    16'd38985: out <= 16'h0516;    16'd38986: out <= 16'h055C;    16'd38987: out <= 16'hFDB7;
    16'd38988: out <= 16'h03B7;    16'd38989: out <= 16'h0158;    16'd38990: out <= 16'h0390;    16'd38991: out <= 16'hFE28;
    16'd38992: out <= 16'h004F;    16'd38993: out <= 16'h005F;    16'd38994: out <= 16'hFF35;    16'd38995: out <= 16'hFB63;
    16'd38996: out <= 16'h06B9;    16'd38997: out <= 16'h0466;    16'd38998: out <= 16'h0512;    16'd38999: out <= 16'hFF40;
    16'd39000: out <= 16'h05E3;    16'd39001: out <= 16'h04FA;    16'd39002: out <= 16'h02B4;    16'd39003: out <= 16'h01C8;
    16'd39004: out <= 16'h0558;    16'd39005: out <= 16'h0A79;    16'd39006: out <= 16'h08CB;    16'd39007: out <= 16'h0240;
    16'd39008: out <= 16'h01C7;    16'd39009: out <= 16'h04AD;    16'd39010: out <= 16'h0B6B;    16'd39011: out <= 16'h039D;
    16'd39012: out <= 16'h052F;    16'd39013: out <= 16'h072B;    16'd39014: out <= 16'h016A;    16'd39015: out <= 16'hFEA0;
    16'd39016: out <= 16'h063D;    16'd39017: out <= 16'h05E4;    16'd39018: out <= 16'h0537;    16'd39019: out <= 16'hFE59;
    16'd39020: out <= 16'h0575;    16'd39021: out <= 16'hFD7A;    16'd39022: out <= 16'h0038;    16'd39023: out <= 16'h0253;
    16'd39024: out <= 16'h0755;    16'd39025: out <= 16'hFEAA;    16'd39026: out <= 16'h0188;    16'd39027: out <= 16'h05FE;
    16'd39028: out <= 16'h035F;    16'd39029: out <= 16'hFDBA;    16'd39030: out <= 16'hFB45;    16'd39031: out <= 16'hFCEB;
    16'd39032: out <= 16'hFD5B;    16'd39033: out <= 16'hFFFB;    16'd39034: out <= 16'hFD7E;    16'd39035: out <= 16'hFFA7;
    16'd39036: out <= 16'h01FC;    16'd39037: out <= 16'h08C9;    16'd39038: out <= 16'h04AB;    16'd39039: out <= 16'hFE67;
    16'd39040: out <= 16'h073A;    16'd39041: out <= 16'h02DD;    16'd39042: out <= 16'h03E9;    16'd39043: out <= 16'h00E9;
    16'd39044: out <= 16'h089B;    16'd39045: out <= 16'h0A3A;    16'd39046: out <= 16'h0670;    16'd39047: out <= 16'h020E;
    16'd39048: out <= 16'h01BA;    16'd39049: out <= 16'h0651;    16'd39050: out <= 16'h0A04;    16'd39051: out <= 16'h0371;
    16'd39052: out <= 16'h07BF;    16'd39053: out <= 16'h0302;    16'd39054: out <= 16'h058F;    16'd39055: out <= 16'hFE6C;
    16'd39056: out <= 16'h0050;    16'd39057: out <= 16'h0265;    16'd39058: out <= 16'h0121;    16'd39059: out <= 16'h02BA;
    16'd39060: out <= 16'h019A;    16'd39061: out <= 16'h02B1;    16'd39062: out <= 16'h008E;    16'd39063: out <= 16'h0495;
    16'd39064: out <= 16'hFFA2;    16'd39065: out <= 16'h03F5;    16'd39066: out <= 16'h0486;    16'd39067: out <= 16'h0226;
    16'd39068: out <= 16'hFE26;    16'd39069: out <= 16'hFD2B;    16'd39070: out <= 16'h0624;    16'd39071: out <= 16'h0675;
    16'd39072: out <= 16'h0233;    16'd39073: out <= 16'h0806;    16'd39074: out <= 16'h04F5;    16'd39075: out <= 16'h002F;
    16'd39076: out <= 16'h03B0;    16'd39077: out <= 16'hF89D;    16'd39078: out <= 16'hFDBA;    16'd39079: out <= 16'h05D1;
    16'd39080: out <= 16'h0441;    16'd39081: out <= 16'hFE8E;    16'd39082: out <= 16'h030A;    16'd39083: out <= 16'h02BA;
    16'd39084: out <= 16'h09C5;    16'd39085: out <= 16'h08C1;    16'd39086: out <= 16'h0154;    16'd39087: out <= 16'h047C;
    16'd39088: out <= 16'h0726;    16'd39089: out <= 16'h00F0;    16'd39090: out <= 16'h00EC;    16'd39091: out <= 16'h0666;
    16'd39092: out <= 16'h0617;    16'd39093: out <= 16'h02AE;    16'd39094: out <= 16'h03AA;    16'd39095: out <= 16'h00CF;
    16'd39096: out <= 16'h054A;    16'd39097: out <= 16'hFDA6;    16'd39098: out <= 16'h0573;    16'd39099: out <= 16'h03F6;
    16'd39100: out <= 16'h07A4;    16'd39101: out <= 16'h05EB;    16'd39102: out <= 16'h05F9;    16'd39103: out <= 16'hFF0E;
    16'd39104: out <= 16'h04B5;    16'd39105: out <= 16'h050A;    16'd39106: out <= 16'h00A8;    16'd39107: out <= 16'h030D;
    16'd39108: out <= 16'h05BD;    16'd39109: out <= 16'h03C3;    16'd39110: out <= 16'h0180;    16'd39111: out <= 16'h07AE;
    16'd39112: out <= 16'h038E;    16'd39113: out <= 16'h0A63;    16'd39114: out <= 16'h0153;    16'd39115: out <= 16'h001F;
    16'd39116: out <= 16'hF775;    16'd39117: out <= 16'h05C3;    16'd39118: out <= 16'h0893;    16'd39119: out <= 16'hF98B;
    16'd39120: out <= 16'h0119;    16'd39121: out <= 16'hFEBE;    16'd39122: out <= 16'hFB20;    16'd39123: out <= 16'h0385;
    16'd39124: out <= 16'hFC18;    16'd39125: out <= 16'hFEA3;    16'd39126: out <= 16'h0388;    16'd39127: out <= 16'hFF4B;
    16'd39128: out <= 16'h08B4;    16'd39129: out <= 16'h01DF;    16'd39130: out <= 16'h03A1;    16'd39131: out <= 16'hFE30;
    16'd39132: out <= 16'h05F1;    16'd39133: out <= 16'hFFDB;    16'd39134: out <= 16'h019F;    16'd39135: out <= 16'h0269;
    16'd39136: out <= 16'h018E;    16'd39137: out <= 16'h043A;    16'd39138: out <= 16'hFFA7;    16'd39139: out <= 16'h075D;
    16'd39140: out <= 16'h069B;    16'd39141: out <= 16'h0408;    16'd39142: out <= 16'h0747;    16'd39143: out <= 16'h0354;
    16'd39144: out <= 16'hFDC3;    16'd39145: out <= 16'h01C0;    16'd39146: out <= 16'hFD25;    16'd39147: out <= 16'h0561;
    16'd39148: out <= 16'h0517;    16'd39149: out <= 16'h03BE;    16'd39150: out <= 16'h0715;    16'd39151: out <= 16'hFC33;
    16'd39152: out <= 16'h0126;    16'd39153: out <= 16'hFAB3;    16'd39154: out <= 16'h036E;    16'd39155: out <= 16'hFBC5;
    16'd39156: out <= 16'hF99C;    16'd39157: out <= 16'h0987;    16'd39158: out <= 16'h002C;    16'd39159: out <= 16'hFD3F;
    16'd39160: out <= 16'h018E;    16'd39161: out <= 16'h0331;    16'd39162: out <= 16'hFF07;    16'd39163: out <= 16'hFDBF;
    16'd39164: out <= 16'h0646;    16'd39165: out <= 16'hFDD9;    16'd39166: out <= 16'hFE94;    16'd39167: out <= 16'h03E3;
    16'd39168: out <= 16'hFD3B;    16'd39169: out <= 16'h00E4;    16'd39170: out <= 16'h03BF;    16'd39171: out <= 16'hF902;
    16'd39172: out <= 16'h00E3;    16'd39173: out <= 16'hFE33;    16'd39174: out <= 16'hF8D9;    16'd39175: out <= 16'hFBAC;
    16'd39176: out <= 16'h0722;    16'd39177: out <= 16'hFF5B;    16'd39178: out <= 16'hFD7D;    16'd39179: out <= 16'h00EF;
    16'd39180: out <= 16'h0286;    16'd39181: out <= 16'h0459;    16'd39182: out <= 16'h00E9;    16'd39183: out <= 16'h0201;
    16'd39184: out <= 16'hFE03;    16'd39185: out <= 16'h0176;    16'd39186: out <= 16'hFD40;    16'd39187: out <= 16'h01DA;
    16'd39188: out <= 16'hFF32;    16'd39189: out <= 16'hFAD3;    16'd39190: out <= 16'hF505;    16'd39191: out <= 16'hFFA0;
    16'd39192: out <= 16'hFE11;    16'd39193: out <= 16'h0267;    16'd39194: out <= 16'hFDF9;    16'd39195: out <= 16'hFCFD;
    16'd39196: out <= 16'hFFD6;    16'd39197: out <= 16'h0960;    16'd39198: out <= 16'h07F2;    16'd39199: out <= 16'hFFB0;
    16'd39200: out <= 16'h0727;    16'd39201: out <= 16'h06B7;    16'd39202: out <= 16'h0513;    16'd39203: out <= 16'h0573;
    16'd39204: out <= 16'h0178;    16'd39205: out <= 16'h0962;    16'd39206: out <= 16'hFF65;    16'd39207: out <= 16'h0162;
    16'd39208: out <= 16'h03AA;    16'd39209: out <= 16'h0304;    16'd39210: out <= 16'h0593;    16'd39211: out <= 16'h0122;
    16'd39212: out <= 16'hFDFD;    16'd39213: out <= 16'h01E4;    16'd39214: out <= 16'h090F;    16'd39215: out <= 16'h0619;
    16'd39216: out <= 16'h022D;    16'd39217: out <= 16'hF9F5;    16'd39218: out <= 16'h026F;    16'd39219: out <= 16'h0407;
    16'd39220: out <= 16'h06F7;    16'd39221: out <= 16'hFB44;    16'd39222: out <= 16'hFCDE;    16'd39223: out <= 16'h06F4;
    16'd39224: out <= 16'h010E;    16'd39225: out <= 16'hFD98;    16'd39226: out <= 16'h0F30;    16'd39227: out <= 16'h06E6;
    16'd39228: out <= 16'h0719;    16'd39229: out <= 16'h062F;    16'd39230: out <= 16'hFD94;    16'd39231: out <= 16'h07B3;
    16'd39232: out <= 16'hFD60;    16'd39233: out <= 16'h0242;    16'd39234: out <= 16'hFD42;    16'd39235: out <= 16'h03F9;
    16'd39236: out <= 16'h0775;    16'd39237: out <= 16'h027F;    16'd39238: out <= 16'h0A9B;    16'd39239: out <= 16'h05F0;
    16'd39240: out <= 16'h0362;    16'd39241: out <= 16'h0195;    16'd39242: out <= 16'h00C3;    16'd39243: out <= 16'h032E;
    16'd39244: out <= 16'h0943;    16'd39245: out <= 16'h05CA;    16'd39246: out <= 16'h0850;    16'd39247: out <= 16'h085E;
    16'd39248: out <= 16'h0494;    16'd39249: out <= 16'h05F7;    16'd39250: out <= 16'h040A;    16'd39251: out <= 16'h01BA;
    16'd39252: out <= 16'h010C;    16'd39253: out <= 16'h00BC;    16'd39254: out <= 16'h008F;    16'd39255: out <= 16'h0499;
    16'd39256: out <= 16'h0133;    16'd39257: out <= 16'h0406;    16'd39258: out <= 16'h0695;    16'd39259: out <= 16'h0D4C;
    16'd39260: out <= 16'h01B7;    16'd39261: out <= 16'h0851;    16'd39262: out <= 16'h05ED;    16'd39263: out <= 16'h0358;
    16'd39264: out <= 16'h017C;    16'd39265: out <= 16'h052C;    16'd39266: out <= 16'hFF27;    16'd39267: out <= 16'h05FE;
    16'd39268: out <= 16'h051A;    16'd39269: out <= 16'hFD6D;    16'd39270: out <= 16'h005E;    16'd39271: out <= 16'h08E9;
    16'd39272: out <= 16'hFED1;    16'd39273: out <= 16'h070D;    16'd39274: out <= 16'h0980;    16'd39275: out <= 16'h043E;
    16'd39276: out <= 16'h050F;    16'd39277: out <= 16'h0807;    16'd39278: out <= 16'h030D;    16'd39279: out <= 16'h0967;
    16'd39280: out <= 16'h02B3;    16'd39281: out <= 16'hFB7C;    16'd39282: out <= 16'hFE35;    16'd39283: out <= 16'h012C;
    16'd39284: out <= 16'hF781;    16'd39285: out <= 16'hFC88;    16'd39286: out <= 16'hFE45;    16'd39287: out <= 16'hF9FA;
    16'd39288: out <= 16'hFE47;    16'd39289: out <= 16'h0954;    16'd39290: out <= 16'h0A8F;    16'd39291: out <= 16'h00FA;
    16'd39292: out <= 16'h05B5;    16'd39293: out <= 16'hFFDB;    16'd39294: out <= 16'h04AD;    16'd39295: out <= 16'h0143;
    16'd39296: out <= 16'h0710;    16'd39297: out <= 16'h0907;    16'd39298: out <= 16'h03F8;    16'd39299: out <= 16'h0922;
    16'd39300: out <= 16'h034F;    16'd39301: out <= 16'h01D4;    16'd39302: out <= 16'h07D4;    16'd39303: out <= 16'h0573;
    16'd39304: out <= 16'h0010;    16'd39305: out <= 16'h01AB;    16'd39306: out <= 16'h0A32;    16'd39307: out <= 16'h02B5;
    16'd39308: out <= 16'h07DE;    16'd39309: out <= 16'h036A;    16'd39310: out <= 16'h03DB;    16'd39311: out <= 16'hFE7F;
    16'd39312: out <= 16'h072D;    16'd39313: out <= 16'hFFBA;    16'd39314: out <= 16'h0492;    16'd39315: out <= 16'hFEEA;
    16'd39316: out <= 16'h06EC;    16'd39317: out <= 16'h035D;    16'd39318: out <= 16'h069D;    16'd39319: out <= 16'h0865;
    16'd39320: out <= 16'h07EF;    16'd39321: out <= 16'h066A;    16'd39322: out <= 16'h01E1;    16'd39323: out <= 16'h0068;
    16'd39324: out <= 16'h0467;    16'd39325: out <= 16'hFF2A;    16'd39326: out <= 16'h00F4;    16'd39327: out <= 16'h06B0;
    16'd39328: out <= 16'h040F;    16'd39329: out <= 16'hFB4B;    16'd39330: out <= 16'h0866;    16'd39331: out <= 16'h0044;
    16'd39332: out <= 16'hFB06;    16'd39333: out <= 16'h0768;    16'd39334: out <= 16'h0218;    16'd39335: out <= 16'h0892;
    16'd39336: out <= 16'h00E9;    16'd39337: out <= 16'h0BB1;    16'd39338: out <= 16'h00E9;    16'd39339: out <= 16'h0816;
    16'd39340: out <= 16'h08D5;    16'd39341: out <= 16'h064A;    16'd39342: out <= 16'h0101;    16'd39343: out <= 16'h00DB;
    16'd39344: out <= 16'h02C2;    16'd39345: out <= 16'h0A29;    16'd39346: out <= 16'hFD89;    16'd39347: out <= 16'h0915;
    16'd39348: out <= 16'h00E7;    16'd39349: out <= 16'h0305;    16'd39350: out <= 16'h0533;    16'd39351: out <= 16'h07BE;
    16'd39352: out <= 16'hFF67;    16'd39353: out <= 16'h05D5;    16'd39354: out <= 16'h0275;    16'd39355: out <= 16'h0813;
    16'd39356: out <= 16'hFF36;    16'd39357: out <= 16'h01AE;    16'd39358: out <= 16'hFD9E;    16'd39359: out <= 16'h070F;
    16'd39360: out <= 16'h0645;    16'd39361: out <= 16'h01D8;    16'd39362: out <= 16'h060C;    16'd39363: out <= 16'hFD09;
    16'd39364: out <= 16'h0395;    16'd39365: out <= 16'h0AA0;    16'd39366: out <= 16'h0452;    16'd39367: out <= 16'h027A;
    16'd39368: out <= 16'h0991;    16'd39369: out <= 16'h024A;    16'd39370: out <= 16'h05ED;    16'd39371: out <= 16'h0139;
    16'd39372: out <= 16'h0631;    16'd39373: out <= 16'hF93A;    16'd39374: out <= 16'h0483;    16'd39375: out <= 16'h0777;
    16'd39376: out <= 16'h010B;    16'd39377: out <= 16'h02D9;    16'd39378: out <= 16'h07F6;    16'd39379: out <= 16'h080D;
    16'd39380: out <= 16'hF92A;    16'd39381: out <= 16'hFE6F;    16'd39382: out <= 16'hFF8D;    16'd39383: out <= 16'h05F0;
    16'd39384: out <= 16'h0562;    16'd39385: out <= 16'h04A8;    16'd39386: out <= 16'hFEA7;    16'd39387: out <= 16'h0221;
    16'd39388: out <= 16'h010A;    16'd39389: out <= 16'h07CB;    16'd39390: out <= 16'h0080;    16'd39391: out <= 16'hFF18;
    16'd39392: out <= 16'h0282;    16'd39393: out <= 16'h0A16;    16'd39394: out <= 16'h090B;    16'd39395: out <= 16'h03B2;
    16'd39396: out <= 16'h0493;    16'd39397: out <= 16'hFFA4;    16'd39398: out <= 16'hFA47;    16'd39399: out <= 16'hFC17;
    16'd39400: out <= 16'hFCE4;    16'd39401: out <= 16'h05A4;    16'd39402: out <= 16'hFD5E;    16'd39403: out <= 16'h061D;
    16'd39404: out <= 16'h00FD;    16'd39405: out <= 16'hFE43;    16'd39406: out <= 16'h0740;    16'd39407: out <= 16'h024F;
    16'd39408: out <= 16'hFCA1;    16'd39409: out <= 16'h02D0;    16'd39410: out <= 16'h01C7;    16'd39411: out <= 16'h03E8;
    16'd39412: out <= 16'h00B3;    16'd39413: out <= 16'h0632;    16'd39414: out <= 16'h0225;    16'd39415: out <= 16'h0AA7;
    16'd39416: out <= 16'h0336;    16'd39417: out <= 16'h01A6;    16'd39418: out <= 16'hFCFC;    16'd39419: out <= 16'h0039;
    16'd39420: out <= 16'h02F9;    16'd39421: out <= 16'h0377;    16'd39422: out <= 16'h0002;    16'd39423: out <= 16'hFFB2;
    16'd39424: out <= 16'h006F;    16'd39425: out <= 16'hFC20;    16'd39426: out <= 16'h03F6;    16'd39427: out <= 16'h01D1;
    16'd39428: out <= 16'hFD17;    16'd39429: out <= 16'hFDE8;    16'd39430: out <= 16'hFF10;    16'd39431: out <= 16'h0667;
    16'd39432: out <= 16'h0612;    16'd39433: out <= 16'hFAEE;    16'd39434: out <= 16'h0031;    16'd39435: out <= 16'h012A;
    16'd39436: out <= 16'hFCDB;    16'd39437: out <= 16'h02F1;    16'd39438: out <= 16'hFF93;    16'd39439: out <= 16'hF827;
    16'd39440: out <= 16'h0455;    16'd39441: out <= 16'h0398;    16'd39442: out <= 16'h0093;    16'd39443: out <= 16'h03D0;
    16'd39444: out <= 16'h07AC;    16'd39445: out <= 16'hFF5E;    16'd39446: out <= 16'h05A7;    16'd39447: out <= 16'hF958;
    16'd39448: out <= 16'h0AE5;    16'd39449: out <= 16'hFB4D;    16'd39450: out <= 16'h01F1;    16'd39451: out <= 16'hFE7F;
    16'd39452: out <= 16'hFF9C;    16'd39453: out <= 16'h00BE;    16'd39454: out <= 16'h02BC;    16'd39455: out <= 16'h0526;
    16'd39456: out <= 16'h0344;    16'd39457: out <= 16'hF9A0;    16'd39458: out <= 16'h02D7;    16'd39459: out <= 16'hFF4E;
    16'd39460: out <= 16'h0350;    16'd39461: out <= 16'h070C;    16'd39462: out <= 16'h0846;    16'd39463: out <= 16'h0E50;
    16'd39464: out <= 16'h051D;    16'd39465: out <= 16'h0A78;    16'd39466: out <= 16'h0449;    16'd39467: out <= 16'h0520;
    16'd39468: out <= 16'h02DD;    16'd39469: out <= 16'h090B;    16'd39470: out <= 16'h06A8;    16'd39471: out <= 16'h06C0;
    16'd39472: out <= 16'h04B5;    16'd39473: out <= 16'h04A9;    16'd39474: out <= 16'h015B;    16'd39475: out <= 16'h0621;
    16'd39476: out <= 16'h00F5;    16'd39477: out <= 16'h02D2;    16'd39478: out <= 16'h05D1;    16'd39479: out <= 16'h025B;
    16'd39480: out <= 16'h03FD;    16'd39481: out <= 16'h046A;    16'd39482: out <= 16'h0689;    16'd39483: out <= 16'h00A3;
    16'd39484: out <= 16'h0495;    16'd39485: out <= 16'h0B44;    16'd39486: out <= 16'h0144;    16'd39487: out <= 16'hFF58;
    16'd39488: out <= 16'h0211;    16'd39489: out <= 16'h052D;    16'd39490: out <= 16'h0417;    16'd39491: out <= 16'h05DE;
    16'd39492: out <= 16'h0452;    16'd39493: out <= 16'h00BD;    16'd39494: out <= 16'h0148;    16'd39495: out <= 16'h034D;
    16'd39496: out <= 16'h039A;    16'd39497: out <= 16'h0487;    16'd39498: out <= 16'hFF16;    16'd39499: out <= 16'hFC65;
    16'd39500: out <= 16'h0641;    16'd39501: out <= 16'h0180;    16'd39502: out <= 16'h0317;    16'd39503: out <= 16'hFD31;
    16'd39504: out <= 16'h025B;    16'd39505: out <= 16'h0710;    16'd39506: out <= 16'h0164;    16'd39507: out <= 16'h0373;
    16'd39508: out <= 16'h0237;    16'd39509: out <= 16'hFF6C;    16'd39510: out <= 16'h00FC;    16'd39511: out <= 16'h0628;
    16'd39512: out <= 16'h03AC;    16'd39513: out <= 16'h04FC;    16'd39514: out <= 16'h05A4;    16'd39515: out <= 16'h065A;
    16'd39516: out <= 16'h0592;    16'd39517: out <= 16'h05B0;    16'd39518: out <= 16'h07A8;    16'd39519: out <= 16'h03FF;
    16'd39520: out <= 16'hFE25;    16'd39521: out <= 16'h0006;    16'd39522: out <= 16'h0745;    16'd39523: out <= 16'h0873;
    16'd39524: out <= 16'h096B;    16'd39525: out <= 16'h0673;    16'd39526: out <= 16'hFF47;    16'd39527: out <= 16'h0722;
    16'd39528: out <= 16'h00C3;    16'd39529: out <= 16'h00C5;    16'd39530: out <= 16'h07B0;    16'd39531: out <= 16'h04C0;
    16'd39532: out <= 16'hFBCA;    16'd39533: out <= 16'hFE34;    16'd39534: out <= 16'h0549;    16'd39535: out <= 16'h0924;
    16'd39536: out <= 16'h04AB;    16'd39537: out <= 16'h022A;    16'd39538: out <= 16'hFDE3;    16'd39539: out <= 16'h010B;
    16'd39540: out <= 16'hFFD5;    16'd39541: out <= 16'hFF0C;    16'd39542: out <= 16'h041C;    16'd39543: out <= 16'hFAD2;
    16'd39544: out <= 16'h01C4;    16'd39545: out <= 16'h07F1;    16'd39546: out <= 16'h02DA;    16'd39547: out <= 16'hFEF8;
    16'd39548: out <= 16'h0525;    16'd39549: out <= 16'h0197;    16'd39550: out <= 16'h03B9;    16'd39551: out <= 16'h03E5;
    16'd39552: out <= 16'h0511;    16'd39553: out <= 16'hFEBC;    16'd39554: out <= 16'h0F87;    16'd39555: out <= 16'h05ED;
    16'd39556: out <= 16'h081E;    16'd39557: out <= 16'h056E;    16'd39558: out <= 16'hFFE7;    16'd39559: out <= 16'h02F0;
    16'd39560: out <= 16'h04C7;    16'd39561: out <= 16'h0181;    16'd39562: out <= 16'h01D4;    16'd39563: out <= 16'h0415;
    16'd39564: out <= 16'hF8F8;    16'd39565: out <= 16'h0046;    16'd39566: out <= 16'h02C8;    16'd39567: out <= 16'h0521;
    16'd39568: out <= 16'h0787;    16'd39569: out <= 16'h0646;    16'd39570: out <= 16'h02A7;    16'd39571: out <= 16'h02E8;
    16'd39572: out <= 16'h0277;    16'd39573: out <= 16'h0851;    16'd39574: out <= 16'h035A;    16'd39575: out <= 16'h0770;
    16'd39576: out <= 16'h02A7;    16'd39577: out <= 16'h0540;    16'd39578: out <= 16'h029F;    16'd39579: out <= 16'hFF3C;
    16'd39580: out <= 16'h02F7;    16'd39581: out <= 16'h0587;    16'd39582: out <= 16'h061E;    16'd39583: out <= 16'h024B;
    16'd39584: out <= 16'h01A9;    16'd39585: out <= 16'h04B3;    16'd39586: out <= 16'h03E4;    16'd39587: out <= 16'h05D2;
    16'd39588: out <= 16'h0707;    16'd39589: out <= 16'h0428;    16'd39590: out <= 16'h0048;    16'd39591: out <= 16'hFECD;
    16'd39592: out <= 16'hFFDB;    16'd39593: out <= 16'hFE21;    16'd39594: out <= 16'h007B;    16'd39595: out <= 16'h0495;
    16'd39596: out <= 16'h04CE;    16'd39597: out <= 16'h04B1;    16'd39598: out <= 16'h06AC;    16'd39599: out <= 16'h037A;
    16'd39600: out <= 16'h0080;    16'd39601: out <= 16'h0553;    16'd39602: out <= 16'hFFF0;    16'd39603: out <= 16'h010D;
    16'd39604: out <= 16'h087C;    16'd39605: out <= 16'h059B;    16'd39606: out <= 16'h018E;    16'd39607: out <= 16'h0062;
    16'd39608: out <= 16'h0898;    16'd39609: out <= 16'h0488;    16'd39610: out <= 16'hFFFB;    16'd39611: out <= 16'h0443;
    16'd39612: out <= 16'h0622;    16'd39613: out <= 16'h079D;    16'd39614: out <= 16'hFDEA;    16'd39615: out <= 16'hFF6A;
    16'd39616: out <= 16'hFDEC;    16'd39617: out <= 16'h0A65;    16'd39618: out <= 16'h00EF;    16'd39619: out <= 16'h0A17;
    16'd39620: out <= 16'hFF04;    16'd39621: out <= 16'h03BA;    16'd39622: out <= 16'h02E8;    16'd39623: out <= 16'h07FB;
    16'd39624: out <= 16'h038A;    16'd39625: out <= 16'h009F;    16'd39626: out <= 16'h0B6A;    16'd39627: out <= 16'h05ED;
    16'd39628: out <= 16'hFCBE;    16'd39629: out <= 16'h09B8;    16'd39630: out <= 16'hFF0F;    16'd39631: out <= 16'hFD9F;
    16'd39632: out <= 16'hFF5C;    16'd39633: out <= 16'h032F;    16'd39634: out <= 16'h001A;    16'd39635: out <= 16'hFDC4;
    16'd39636: out <= 16'h03BD;    16'd39637: out <= 16'h034B;    16'd39638: out <= 16'h0613;    16'd39639: out <= 16'h064E;
    16'd39640: out <= 16'hFD54;    16'd39641: out <= 16'hFE08;    16'd39642: out <= 16'h05DB;    16'd39643: out <= 16'h04E3;
    16'd39644: out <= 16'h01C9;    16'd39645: out <= 16'h00CC;    16'd39646: out <= 16'h0BB4;    16'd39647: out <= 16'h06BE;
    16'd39648: out <= 16'h018E;    16'd39649: out <= 16'h0118;    16'd39650: out <= 16'h0357;    16'd39651: out <= 16'h00E5;
    16'd39652: out <= 16'h038C;    16'd39653: out <= 16'h0184;    16'd39654: out <= 16'h0421;    16'd39655: out <= 16'hFE39;
    16'd39656: out <= 16'hFC8F;    16'd39657: out <= 16'h051D;    16'd39658: out <= 16'h01E4;    16'd39659: out <= 16'h04D7;
    16'd39660: out <= 16'hFA79;    16'd39661: out <= 16'h075D;    16'd39662: out <= 16'h0253;    16'd39663: out <= 16'h069D;
    16'd39664: out <= 16'h03CC;    16'd39665: out <= 16'hFCC3;    16'd39666: out <= 16'hFDAD;    16'd39667: out <= 16'h02B5;
    16'd39668: out <= 16'h00CA;    16'd39669: out <= 16'h02F4;    16'd39670: out <= 16'hFFE3;    16'd39671: out <= 16'h03A6;
    16'd39672: out <= 16'hFAEF;    16'd39673: out <= 16'h0131;    16'd39674: out <= 16'h01B4;    16'd39675: out <= 16'hFACA;
    16'd39676: out <= 16'h00DA;    16'd39677: out <= 16'hFEEC;    16'd39678: out <= 16'hFF95;    16'd39679: out <= 16'h0568;
    16'd39680: out <= 16'h08C4;    16'd39681: out <= 16'h01C3;    16'd39682: out <= 16'hFB46;    16'd39683: out <= 16'hFF18;
    16'd39684: out <= 16'h0144;    16'd39685: out <= 16'h021A;    16'd39686: out <= 16'hF824;    16'd39687: out <= 16'hFF58;
    16'd39688: out <= 16'h012D;    16'd39689: out <= 16'hFD05;    16'd39690: out <= 16'hFE5E;    16'd39691: out <= 16'h03CE;
    16'd39692: out <= 16'h0356;    16'd39693: out <= 16'hFD1E;    16'd39694: out <= 16'hFB65;    16'd39695: out <= 16'h0319;
    16'd39696: out <= 16'hFBA0;    16'd39697: out <= 16'hF9B7;    16'd39698: out <= 16'hFDCB;    16'd39699: out <= 16'hFCF3;
    16'd39700: out <= 16'hFD6F;    16'd39701: out <= 16'h04E4;    16'd39702: out <= 16'hFFD0;    16'd39703: out <= 16'hFF9F;
    16'd39704: out <= 16'hFA9B;    16'd39705: out <= 16'hFDE1;    16'd39706: out <= 16'h045A;    16'd39707: out <= 16'hFF5B;
    16'd39708: out <= 16'hFD9B;    16'd39709: out <= 16'h013F;    16'd39710: out <= 16'h01FB;    16'd39711: out <= 16'h02F2;
    16'd39712: out <= 16'h00C6;    16'd39713: out <= 16'h009C;    16'd39714: out <= 16'h02A3;    16'd39715: out <= 16'h0220;
    16'd39716: out <= 16'h06E1;    16'd39717: out <= 16'h0764;    16'd39718: out <= 16'h0561;    16'd39719: out <= 16'h0455;
    16'd39720: out <= 16'h01FB;    16'd39721: out <= 16'h0B10;    16'd39722: out <= 16'h0261;    16'd39723: out <= 16'h063E;
    16'd39724: out <= 16'h0782;    16'd39725: out <= 16'h0794;    16'd39726: out <= 16'h023A;    16'd39727: out <= 16'h0A32;
    16'd39728: out <= 16'h08AB;    16'd39729: out <= 16'h08DD;    16'd39730: out <= 16'h01FC;    16'd39731: out <= 16'h00C2;
    16'd39732: out <= 16'h017D;    16'd39733: out <= 16'h0100;    16'd39734: out <= 16'h0253;    16'd39735: out <= 16'h0524;
    16'd39736: out <= 16'h01A8;    16'd39737: out <= 16'h079E;    16'd39738: out <= 16'h01D0;    16'd39739: out <= 16'hFFC1;
    16'd39740: out <= 16'h081F;    16'd39741: out <= 16'h06CC;    16'd39742: out <= 16'h0736;    16'd39743: out <= 16'h0471;
    16'd39744: out <= 16'h08E6;    16'd39745: out <= 16'h06DA;    16'd39746: out <= 16'h06F2;    16'd39747: out <= 16'h012A;
    16'd39748: out <= 16'h022D;    16'd39749: out <= 16'h0678;    16'd39750: out <= 16'h0220;    16'd39751: out <= 16'h0C57;
    16'd39752: out <= 16'h070C;    16'd39753: out <= 16'h0989;    16'd39754: out <= 16'hFBE4;    16'd39755: out <= 16'h0129;
    16'd39756: out <= 16'h0500;    16'd39757: out <= 16'h04EA;    16'd39758: out <= 16'hFF13;    16'd39759: out <= 16'h010C;
    16'd39760: out <= 16'h0665;    16'd39761: out <= 16'h0A46;    16'd39762: out <= 16'h026E;    16'd39763: out <= 16'h072E;
    16'd39764: out <= 16'h0261;    16'd39765: out <= 16'h04B2;    16'd39766: out <= 16'h04C6;    16'd39767: out <= 16'hFE57;
    16'd39768: out <= 16'h03E8;    16'd39769: out <= 16'h0151;    16'd39770: out <= 16'h07EC;    16'd39771: out <= 16'h08E7;
    16'd39772: out <= 16'h01C2;    16'd39773: out <= 16'hFFD5;    16'd39774: out <= 16'h0655;    16'd39775: out <= 16'h08D6;
    16'd39776: out <= 16'hFFD1;    16'd39777: out <= 16'h0050;    16'd39778: out <= 16'h009C;    16'd39779: out <= 16'h06FF;
    16'd39780: out <= 16'h05E7;    16'd39781: out <= 16'hFFD6;    16'd39782: out <= 16'h029E;    16'd39783: out <= 16'hFD52;
    16'd39784: out <= 16'h0AC1;    16'd39785: out <= 16'h0D77;    16'd39786: out <= 16'h013A;    16'd39787: out <= 16'h05E0;
    16'd39788: out <= 16'h0562;    16'd39789: out <= 16'h03A1;    16'd39790: out <= 16'h07CB;    16'd39791: out <= 16'hFF19;
    16'd39792: out <= 16'h037A;    16'd39793: out <= 16'h0130;    16'd39794: out <= 16'h06EF;    16'd39795: out <= 16'h00B3;
    16'd39796: out <= 16'hFC10;    16'd39797: out <= 16'h0268;    16'd39798: out <= 16'h0516;    16'd39799: out <= 16'hF9C5;
    16'd39800: out <= 16'h08BD;    16'd39801: out <= 16'h01AB;    16'd39802: out <= 16'h03FC;    16'd39803: out <= 16'h0A3C;
    16'd39804: out <= 16'h0032;    16'd39805: out <= 16'h0AD7;    16'd39806: out <= 16'h075A;    16'd39807: out <= 16'h05B1;
    16'd39808: out <= 16'h0724;    16'd39809: out <= 16'h035B;    16'd39810: out <= 16'h07D1;    16'd39811: out <= 16'h08DE;
    16'd39812: out <= 16'h07E4;    16'd39813: out <= 16'h0433;    16'd39814: out <= 16'hFF03;    16'd39815: out <= 16'h0159;
    16'd39816: out <= 16'h029C;    16'd39817: out <= 16'h0382;    16'd39818: out <= 16'h0C0C;    16'd39819: out <= 16'hFF5C;
    16'd39820: out <= 16'h01D6;    16'd39821: out <= 16'h0499;    16'd39822: out <= 16'h02FA;    16'd39823: out <= 16'h05AE;
    16'd39824: out <= 16'hFFB8;    16'd39825: out <= 16'h0498;    16'd39826: out <= 16'h07B5;    16'd39827: out <= 16'h0199;
    16'd39828: out <= 16'hFF3B;    16'd39829: out <= 16'h0881;    16'd39830: out <= 16'h00B4;    16'd39831: out <= 16'h0079;
    16'd39832: out <= 16'h049C;    16'd39833: out <= 16'h0578;    16'd39834: out <= 16'h0959;    16'd39835: out <= 16'h0546;
    16'd39836: out <= 16'h0311;    16'd39837: out <= 16'h07BC;    16'd39838: out <= 16'h0550;    16'd39839: out <= 16'h01A4;
    16'd39840: out <= 16'h0801;    16'd39841: out <= 16'h0B35;    16'd39842: out <= 16'h0653;    16'd39843: out <= 16'h0629;
    16'd39844: out <= 16'h042F;    16'd39845: out <= 16'h00E5;    16'd39846: out <= 16'hFE38;    16'd39847: out <= 16'h040F;
    16'd39848: out <= 16'hFEA8;    16'd39849: out <= 16'h0068;    16'd39850: out <= 16'hFFB3;    16'd39851: out <= 16'hFDB5;
    16'd39852: out <= 16'h0522;    16'd39853: out <= 16'h098B;    16'd39854: out <= 16'h018B;    16'd39855: out <= 16'h07D5;
    16'd39856: out <= 16'h0572;    16'd39857: out <= 16'h064D;    16'd39858: out <= 16'h0409;    16'd39859: out <= 16'h043C;
    16'd39860: out <= 16'h0860;    16'd39861: out <= 16'h043A;    16'd39862: out <= 16'h015E;    16'd39863: out <= 16'h0C51;
    16'd39864: out <= 16'h01DA;    16'd39865: out <= 16'h04F4;    16'd39866: out <= 16'h05DD;    16'd39867: out <= 16'h0419;
    16'd39868: out <= 16'h0846;    16'd39869: out <= 16'h0088;    16'd39870: out <= 16'h0238;    16'd39871: out <= 16'h0704;
    16'd39872: out <= 16'h03F0;    16'd39873: out <= 16'h0ADD;    16'd39874: out <= 16'h09EE;    16'd39875: out <= 16'hFFE6;
    16'd39876: out <= 16'hFE42;    16'd39877: out <= 16'h01DB;    16'd39878: out <= 16'h0303;    16'd39879: out <= 16'h03E0;
    16'd39880: out <= 16'h0187;    16'd39881: out <= 16'hF8CC;    16'd39882: out <= 16'h01DE;    16'd39883: out <= 16'h02C7;
    16'd39884: out <= 16'h070F;    16'd39885: out <= 16'h0356;    16'd39886: out <= 16'h0791;    16'd39887: out <= 16'h098F;
    16'd39888: out <= 16'h07FE;    16'd39889: out <= 16'h00B0;    16'd39890: out <= 16'hFF52;    16'd39891: out <= 16'hFEF5;
    16'd39892: out <= 16'h05EC;    16'd39893: out <= 16'h05E9;    16'd39894: out <= 16'h060E;    16'd39895: out <= 16'h0C15;
    16'd39896: out <= 16'h00B8;    16'd39897: out <= 16'h0329;    16'd39898: out <= 16'h0AF8;    16'd39899: out <= 16'h089C;
    16'd39900: out <= 16'h002E;    16'd39901: out <= 16'h0223;    16'd39902: out <= 16'h045B;    16'd39903: out <= 16'hFEEF;
    16'd39904: out <= 16'h0109;    16'd39905: out <= 16'h025F;    16'd39906: out <= 16'h00D6;    16'd39907: out <= 16'h06DE;
    16'd39908: out <= 16'h03C8;    16'd39909: out <= 16'hFE41;    16'd39910: out <= 16'h033E;    16'd39911: out <= 16'h0089;
    16'd39912: out <= 16'h0605;    16'd39913: out <= 16'h0A84;    16'd39914: out <= 16'h01AD;    16'd39915: out <= 16'h0555;
    16'd39916: out <= 16'h0598;    16'd39917: out <= 16'hF936;    16'd39918: out <= 16'hFD0B;    16'd39919: out <= 16'h0063;
    16'd39920: out <= 16'h0605;    16'd39921: out <= 16'hFD83;    16'd39922: out <= 16'h0200;    16'd39923: out <= 16'h0663;
    16'd39924: out <= 16'h06B6;    16'd39925: out <= 16'hFD3A;    16'd39926: out <= 16'h00D5;    16'd39927: out <= 16'h0163;
    16'd39928: out <= 16'h01D1;    16'd39929: out <= 16'h051D;    16'd39930: out <= 16'hFF42;    16'd39931: out <= 16'h04A0;
    16'd39932: out <= 16'h03D2;    16'd39933: out <= 16'hF9A0;    16'd39934: out <= 16'hFE33;    16'd39935: out <= 16'hFC96;
    16'd39936: out <= 16'hFE9D;    16'd39937: out <= 16'hFAF6;    16'd39938: out <= 16'hFE0A;    16'd39939: out <= 16'h0187;
    16'd39940: out <= 16'hFEC3;    16'd39941: out <= 16'h01FE;    16'd39942: out <= 16'hFDE6;    16'd39943: out <= 16'hFBAF;
    16'd39944: out <= 16'h08B3;    16'd39945: out <= 16'h0363;    16'd39946: out <= 16'h050A;    16'd39947: out <= 16'hF5B7;
    16'd39948: out <= 16'h0381;    16'd39949: out <= 16'hFE7F;    16'd39950: out <= 16'h0090;    16'd39951: out <= 16'hFA73;
    16'd39952: out <= 16'hFB3D;    16'd39953: out <= 16'hFF8F;    16'd39954: out <= 16'h00D2;    16'd39955: out <= 16'h05B0;
    16'd39956: out <= 16'h01BA;    16'd39957: out <= 16'hFF42;    16'd39958: out <= 16'hFD92;    16'd39959: out <= 16'hFF7C;
    16'd39960: out <= 16'h02CE;    16'd39961: out <= 16'h033E;    16'd39962: out <= 16'hFAA8;    16'd39963: out <= 16'h031C;
    16'd39964: out <= 16'h0003;    16'd39965: out <= 16'hF907;    16'd39966: out <= 16'h024B;    16'd39967: out <= 16'h05A6;
    16'd39968: out <= 16'hFDFF;    16'd39969: out <= 16'h034C;    16'd39970: out <= 16'h0063;    16'd39971: out <= 16'h0485;
    16'd39972: out <= 16'h048A;    16'd39973: out <= 16'h057E;    16'd39974: out <= 16'hFED4;    16'd39975: out <= 16'h09EC;
    16'd39976: out <= 16'h0732;    16'd39977: out <= 16'h060F;    16'd39978: out <= 16'h06A5;    16'd39979: out <= 16'h0193;
    16'd39980: out <= 16'h0252;    16'd39981: out <= 16'h0155;    16'd39982: out <= 16'hFEEA;    16'd39983: out <= 16'hFFE5;
    16'd39984: out <= 16'h0542;    16'd39985: out <= 16'h032D;    16'd39986: out <= 16'h03B1;    16'd39987: out <= 16'h06BB;
    16'd39988: out <= 16'h084B;    16'd39989: out <= 16'h02EF;    16'd39990: out <= 16'h022F;    16'd39991: out <= 16'h0514;
    16'd39992: out <= 16'h06A7;    16'd39993: out <= 16'hFFC1;    16'd39994: out <= 16'h03D1;    16'd39995: out <= 16'h02CD;
    16'd39996: out <= 16'hFFDD;    16'd39997: out <= 16'h0148;    16'd39998: out <= 16'h01FD;    16'd39999: out <= 16'hFDDC;
    16'd40000: out <= 16'h017C;    16'd40001: out <= 16'hFDBB;    16'd40002: out <= 16'h058B;    16'd40003: out <= 16'hFE74;
    16'd40004: out <= 16'h0051;    16'd40005: out <= 16'h0710;    16'd40006: out <= 16'h0691;    16'd40007: out <= 16'h0879;
    16'd40008: out <= 16'hFD7E;    16'd40009: out <= 16'h0802;    16'd40010: out <= 16'h042B;    16'd40011: out <= 16'hFF24;
    16'd40012: out <= 16'h02FB;    16'd40013: out <= 16'h0671;    16'd40014: out <= 16'h00F4;    16'd40015: out <= 16'h032C;
    16'd40016: out <= 16'h051F;    16'd40017: out <= 16'h0C34;    16'd40018: out <= 16'h0DC3;    16'd40019: out <= 16'h06D8;
    16'd40020: out <= 16'h089C;    16'd40021: out <= 16'h0ADF;    16'd40022: out <= 16'h08B0;    16'd40023: out <= 16'h062A;
    16'd40024: out <= 16'h05E0;    16'd40025: out <= 16'h0A94;    16'd40026: out <= 16'h00B7;    16'd40027: out <= 16'h07FC;
    16'd40028: out <= 16'h0165;    16'd40029: out <= 16'h064C;    16'd40030: out <= 16'h00FE;    16'd40031: out <= 16'h0612;
    16'd40032: out <= 16'h03A7;    16'd40033: out <= 16'h051C;    16'd40034: out <= 16'hFF1B;    16'd40035: out <= 16'h005A;
    16'd40036: out <= 16'h0419;    16'd40037: out <= 16'h041E;    16'd40038: out <= 16'h01E5;    16'd40039: out <= 16'h0032;
    16'd40040: out <= 16'h0417;    16'd40041: out <= 16'h04AA;    16'd40042: out <= 16'h0773;    16'd40043: out <= 16'h0799;
    16'd40044: out <= 16'h03F1;    16'd40045: out <= 16'h076A;    16'd40046: out <= 16'h090B;    16'd40047: out <= 16'h01F6;
    16'd40048: out <= 16'h03AF;    16'd40049: out <= 16'hFC24;    16'd40050: out <= 16'h0014;    16'd40051: out <= 16'hFFBB;
    16'd40052: out <= 16'hFCDF;    16'd40053: out <= 16'hF7D9;    16'd40054: out <= 16'h04FD;    16'd40055: out <= 16'hFF63;
    16'd40056: out <= 16'hFD8B;    16'd40057: out <= 16'hFEB1;    16'd40058: out <= 16'hFF5D;    16'd40059: out <= 16'hFF70;
    16'd40060: out <= 16'h0661;    16'd40061: out <= 16'h0C15;    16'd40062: out <= 16'hFF23;    16'd40063: out <= 16'hFD6B;
    16'd40064: out <= 16'h0518;    16'd40065: out <= 16'h082C;    16'd40066: out <= 16'h0216;    16'd40067: out <= 16'h017B;
    16'd40068: out <= 16'h03E3;    16'd40069: out <= 16'hFF49;    16'd40070: out <= 16'h0312;    16'd40071: out <= 16'hFE83;
    16'd40072: out <= 16'h0161;    16'd40073: out <= 16'h00DD;    16'd40074: out <= 16'hF831;    16'd40075: out <= 16'h0291;
    16'd40076: out <= 16'h04C1;    16'd40077: out <= 16'h06C2;    16'd40078: out <= 16'h01BA;    16'd40079: out <= 16'h068F;
    16'd40080: out <= 16'h02F9;    16'd40081: out <= 16'h051D;    16'd40082: out <= 16'h0000;    16'd40083: out <= 16'h0DA9;
    16'd40084: out <= 16'h005E;    16'd40085: out <= 16'h03D0;    16'd40086: out <= 16'h02A2;    16'd40087: out <= 16'h0305;
    16'd40088: out <= 16'hFE44;    16'd40089: out <= 16'h066A;    16'd40090: out <= 16'hF920;    16'd40091: out <= 16'h009F;
    16'd40092: out <= 16'h0B99;    16'd40093: out <= 16'h06D3;    16'd40094: out <= 16'h0281;    16'd40095: out <= 16'h027A;
    16'd40096: out <= 16'h0145;    16'd40097: out <= 16'h03E2;    16'd40098: out <= 16'h079F;    16'd40099: out <= 16'hFE8A;
    16'd40100: out <= 16'h09A5;    16'd40101: out <= 16'h06F4;    16'd40102: out <= 16'hFEE1;    16'd40103: out <= 16'h03CF;
    16'd40104: out <= 16'h0590;    16'd40105: out <= 16'h022D;    16'd40106: out <= 16'h0250;    16'd40107: out <= 16'h022F;
    16'd40108: out <= 16'hFD39;    16'd40109: out <= 16'h03FE;    16'd40110: out <= 16'h06E9;    16'd40111: out <= 16'h04FF;
    16'd40112: out <= 16'hFF0B;    16'd40113: out <= 16'h0237;    16'd40114: out <= 16'h07B2;    16'd40115: out <= 16'h05A4;
    16'd40116: out <= 16'h03C8;    16'd40117: out <= 16'h0193;    16'd40118: out <= 16'h0270;    16'd40119: out <= 16'h0574;
    16'd40120: out <= 16'h02A2;    16'd40121: out <= 16'h072F;    16'd40122: out <= 16'h01E0;    16'd40123: out <= 16'h01C1;
    16'd40124: out <= 16'h06AB;    16'd40125: out <= 16'h0B0F;    16'd40126: out <= 16'h062D;    16'd40127: out <= 16'h0AC3;
    16'd40128: out <= 16'h0138;    16'd40129: out <= 16'h0652;    16'd40130: out <= 16'h0B9A;    16'd40131: out <= 16'h03A8;
    16'd40132: out <= 16'h0692;    16'd40133: out <= 16'h0901;    16'd40134: out <= 16'h068E;    16'd40135: out <= 16'h06D6;
    16'd40136: out <= 16'h007C;    16'd40137: out <= 16'h0798;    16'd40138: out <= 16'h029D;    16'd40139: out <= 16'h0576;
    16'd40140: out <= 16'h00F1;    16'd40141: out <= 16'h01E1;    16'd40142: out <= 16'h0383;    16'd40143: out <= 16'h0265;
    16'd40144: out <= 16'h00A3;    16'd40145: out <= 16'h06AF;    16'd40146: out <= 16'h0779;    16'd40147: out <= 16'h0133;
    16'd40148: out <= 16'hFCE4;    16'd40149: out <= 16'h035C;    16'd40150: out <= 16'h0625;    16'd40151: out <= 16'h06E1;
    16'd40152: out <= 16'h0156;    16'd40153: out <= 16'h09CC;    16'd40154: out <= 16'h039E;    16'd40155: out <= 16'h0838;
    16'd40156: out <= 16'h042D;    16'd40157: out <= 16'h0268;    16'd40158: out <= 16'h014A;    16'd40159: out <= 16'h03F1;
    16'd40160: out <= 16'hFEF3;    16'd40161: out <= 16'h0335;    16'd40162: out <= 16'h0322;    16'd40163: out <= 16'h00A1;
    16'd40164: out <= 16'h0751;    16'd40165: out <= 16'h02DD;    16'd40166: out <= 16'h0108;    16'd40167: out <= 16'h00C0;
    16'd40168: out <= 16'hFFA8;    16'd40169: out <= 16'h01A7;    16'd40170: out <= 16'h0443;    16'd40171: out <= 16'h06BB;
    16'd40172: out <= 16'hFF60;    16'd40173: out <= 16'h04CF;    16'd40174: out <= 16'h009D;    16'd40175: out <= 16'h0108;
    16'd40176: out <= 16'hFD05;    16'd40177: out <= 16'hFB53;    16'd40178: out <= 16'h06B4;    16'd40179: out <= 16'hFC6E;
    16'd40180: out <= 16'h05F8;    16'd40181: out <= 16'hFC2F;    16'd40182: out <= 16'hFE9F;    16'd40183: out <= 16'hFB36;
    16'd40184: out <= 16'h0202;    16'd40185: out <= 16'hF8C8;    16'd40186: out <= 16'hFDF9;    16'd40187: out <= 16'h071F;
    16'd40188: out <= 16'hFBD8;    16'd40189: out <= 16'hF84D;    16'd40190: out <= 16'h01CB;    16'd40191: out <= 16'h009D;
    16'd40192: out <= 16'hFE93;    16'd40193: out <= 16'h00A9;    16'd40194: out <= 16'h0217;    16'd40195: out <= 16'h0106;
    16'd40196: out <= 16'h02E8;    16'd40197: out <= 16'h016C;    16'd40198: out <= 16'h092B;    16'd40199: out <= 16'hFFF5;
    16'd40200: out <= 16'hFF16;    16'd40201: out <= 16'hFF9E;    16'd40202: out <= 16'hFD95;    16'd40203: out <= 16'h0883;
    16'd40204: out <= 16'hFE32;    16'd40205: out <= 16'h054F;    16'd40206: out <= 16'hFE55;    16'd40207: out <= 16'h0091;
    16'd40208: out <= 16'hF841;    16'd40209: out <= 16'hFCB6;    16'd40210: out <= 16'h0659;    16'd40211: out <= 16'hFEC5;
    16'd40212: out <= 16'h06A1;    16'd40213: out <= 16'h0357;    16'd40214: out <= 16'h022A;    16'd40215: out <= 16'h00B4;
    16'd40216: out <= 16'hFF08;    16'd40217: out <= 16'hFEAC;    16'd40218: out <= 16'hFD61;    16'd40219: out <= 16'hF990;
    16'd40220: out <= 16'hFB14;    16'd40221: out <= 16'h0650;    16'd40222: out <= 16'h0A48;    16'd40223: out <= 16'h045D;
    16'd40224: out <= 16'h0017;    16'd40225: out <= 16'h073D;    16'd40226: out <= 16'hFF5F;    16'd40227: out <= 16'hF9CF;
    16'd40228: out <= 16'h03E2;    16'd40229: out <= 16'h02D8;    16'd40230: out <= 16'h0698;    16'd40231: out <= 16'h0DFB;
    16'd40232: out <= 16'h0604;    16'd40233: out <= 16'h0D45;    16'd40234: out <= 16'h0351;    16'd40235: out <= 16'hFF17;
    16'd40236: out <= 16'h010C;    16'd40237: out <= 16'h0836;    16'd40238: out <= 16'h03D4;    16'd40239: out <= 16'h0091;
    16'd40240: out <= 16'h014F;    16'd40241: out <= 16'h0359;    16'd40242: out <= 16'h034E;    16'd40243: out <= 16'h00F6;
    16'd40244: out <= 16'h0469;    16'd40245: out <= 16'hFD0A;    16'd40246: out <= 16'h078A;    16'd40247: out <= 16'h02E0;
    16'd40248: out <= 16'h03E9;    16'd40249: out <= 16'h0842;    16'd40250: out <= 16'h00BF;    16'd40251: out <= 16'h06A0;
    16'd40252: out <= 16'h07AE;    16'd40253: out <= 16'h035D;    16'd40254: out <= 16'hFD7B;    16'd40255: out <= 16'h08A6;
    16'd40256: out <= 16'h09F6;    16'd40257: out <= 16'h0772;    16'd40258: out <= 16'h03DF;    16'd40259: out <= 16'h017A;
    16'd40260: out <= 16'h0338;    16'd40261: out <= 16'h0D69;    16'd40262: out <= 16'h03A8;    16'd40263: out <= 16'h0913;
    16'd40264: out <= 16'h0B0A;    16'd40265: out <= 16'h02E3;    16'd40266: out <= 16'h03A8;    16'd40267: out <= 16'hFBD0;
    16'd40268: out <= 16'h02CD;    16'd40269: out <= 16'h01DD;    16'd40270: out <= 16'h022B;    16'd40271: out <= 16'h012B;
    16'd40272: out <= 16'h017D;    16'd40273: out <= 16'h038D;    16'd40274: out <= 16'h05A3;    16'd40275: out <= 16'h0278;
    16'd40276: out <= 16'h0627;    16'd40277: out <= 16'h025D;    16'd40278: out <= 16'hFE47;    16'd40279: out <= 16'hFFFD;
    16'd40280: out <= 16'h09A3;    16'd40281: out <= 16'h0372;    16'd40282: out <= 16'h065C;    16'd40283: out <= 16'hFE27;
    16'd40284: out <= 16'h00ED;    16'd40285: out <= 16'h03B9;    16'd40286: out <= 16'h06EE;    16'd40287: out <= 16'h0182;
    16'd40288: out <= 16'h0054;    16'd40289: out <= 16'h0031;    16'd40290: out <= 16'h0419;    16'd40291: out <= 16'hFFF3;
    16'd40292: out <= 16'h03F6;    16'd40293: out <= 16'hFEC1;    16'd40294: out <= 16'h0072;    16'd40295: out <= 16'h0043;
    16'd40296: out <= 16'h025B;    16'd40297: out <= 16'h0742;    16'd40298: out <= 16'h043D;    16'd40299: out <= 16'h0A18;
    16'd40300: out <= 16'h0386;    16'd40301: out <= 16'h068B;    16'd40302: out <= 16'hFFDE;    16'd40303: out <= 16'hF9DF;
    16'd40304: out <= 16'hFF58;    16'd40305: out <= 16'h01D7;    16'd40306: out <= 16'hFDF9;    16'd40307: out <= 16'h00D9;
    16'd40308: out <= 16'h03CD;    16'd40309: out <= 16'hFFCB;    16'd40310: out <= 16'h030E;    16'd40311: out <= 16'h084F;
    16'd40312: out <= 16'hFF21;    16'd40313: out <= 16'h075C;    16'd40314: out <= 16'h08AD;    16'd40315: out <= 16'h04BC;
    16'd40316: out <= 16'hFF77;    16'd40317: out <= 16'h0288;    16'd40318: out <= 16'h0A87;    16'd40319: out <= 16'h0AB2;
    16'd40320: out <= 16'hFCC1;    16'd40321: out <= 16'h06B7;    16'd40322: out <= 16'h02D0;    16'd40323: out <= 16'h089F;
    16'd40324: out <= 16'h02EB;    16'd40325: out <= 16'h058D;    16'd40326: out <= 16'h07CD;    16'd40327: out <= 16'h01F3;
    16'd40328: out <= 16'h046E;    16'd40329: out <= 16'h077B;    16'd40330: out <= 16'h0209;    16'd40331: out <= 16'hFE8C;
    16'd40332: out <= 16'h01B8;    16'd40333: out <= 16'h01B5;    16'd40334: out <= 16'h05BD;    16'd40335: out <= 16'h03F0;
    16'd40336: out <= 16'h0B8C;    16'd40337: out <= 16'h0112;    16'd40338: out <= 16'h0770;    16'd40339: out <= 16'h09C4;
    16'd40340: out <= 16'h033C;    16'd40341: out <= 16'h042A;    16'd40342: out <= 16'h0394;    16'd40343: out <= 16'hFF0F;
    16'd40344: out <= 16'hFF77;    16'd40345: out <= 16'h03C1;    16'd40346: out <= 16'h0393;    16'd40347: out <= 16'h0647;
    16'd40348: out <= 16'hFE25;    16'd40349: out <= 16'h065D;    16'd40350: out <= 16'h02B4;    16'd40351: out <= 16'h027F;
    16'd40352: out <= 16'h037E;    16'd40353: out <= 16'h0231;    16'd40354: out <= 16'h02EA;    16'd40355: out <= 16'hFF5C;
    16'd40356: out <= 16'h08F6;    16'd40357: out <= 16'h0180;    16'd40358: out <= 16'hFDA9;    16'd40359: out <= 16'h0209;
    16'd40360: out <= 16'h09A5;    16'd40361: out <= 16'h0644;    16'd40362: out <= 16'h00D0;    16'd40363: out <= 16'h0541;
    16'd40364: out <= 16'hFD4B;    16'd40365: out <= 16'h0524;    16'd40366: out <= 16'h09D2;    16'd40367: out <= 16'h098C;
    16'd40368: out <= 16'h0541;    16'd40369: out <= 16'h03CF;    16'd40370: out <= 16'h046F;    16'd40371: out <= 16'h0687;
    16'd40372: out <= 16'hFE3E;    16'd40373: out <= 16'h08FD;    16'd40374: out <= 16'h00F8;    16'd40375: out <= 16'h014C;
    16'd40376: out <= 16'h0291;    16'd40377: out <= 16'h0721;    16'd40378: out <= 16'h0B63;    16'd40379: out <= 16'hFFF8;
    16'd40380: out <= 16'h02A8;    16'd40381: out <= 16'h04B3;    16'd40382: out <= 16'h02A7;    16'd40383: out <= 16'h0277;
    16'd40384: out <= 16'h02E0;    16'd40385: out <= 16'h01C4;    16'd40386: out <= 16'h09C0;    16'd40387: out <= 16'h02B6;
    16'd40388: out <= 16'h021A;    16'd40389: out <= 16'h025E;    16'd40390: out <= 16'h065E;    16'd40391: out <= 16'h011F;
    16'd40392: out <= 16'h01C5;    16'd40393: out <= 16'h0497;    16'd40394: out <= 16'h06A5;    16'd40395: out <= 16'h01B8;
    16'd40396: out <= 16'hFE86;    16'd40397: out <= 16'h0196;    16'd40398: out <= 16'h04A3;    16'd40399: out <= 16'h0413;
    16'd40400: out <= 16'h018E;    16'd40401: out <= 16'h05B5;    16'd40402: out <= 16'h056E;    16'd40403: out <= 16'h053E;
    16'd40404: out <= 16'h0275;    16'd40405: out <= 16'h0675;    16'd40406: out <= 16'h0AAE;    16'd40407: out <= 16'hFF42;
    16'd40408: out <= 16'h0231;    16'd40409: out <= 16'hFD66;    16'd40410: out <= 16'h0680;    16'd40411: out <= 16'h01AA;
    16'd40412: out <= 16'h07C8;    16'd40413: out <= 16'h05AD;    16'd40414: out <= 16'h0558;    16'd40415: out <= 16'h03B4;
    16'd40416: out <= 16'h0A0D;    16'd40417: out <= 16'h0645;    16'd40418: out <= 16'h0770;    16'd40419: out <= 16'h0089;
    16'd40420: out <= 16'h0723;    16'd40421: out <= 16'hFF90;    16'd40422: out <= 16'hFBBF;    16'd40423: out <= 16'hFC74;
    16'd40424: out <= 16'hFF00;    16'd40425: out <= 16'hFDE4;    16'd40426: out <= 16'h0548;    16'd40427: out <= 16'hFBF5;
    16'd40428: out <= 16'hFAA3;    16'd40429: out <= 16'h0093;    16'd40430: out <= 16'hF477;    16'd40431: out <= 16'hFD35;
    16'd40432: out <= 16'h022E;    16'd40433: out <= 16'h02C5;    16'd40434: out <= 16'h0176;    16'd40435: out <= 16'hFF44;
    16'd40436: out <= 16'h00D4;    16'd40437: out <= 16'hFBFA;    16'd40438: out <= 16'h05A9;    16'd40439: out <= 16'hF9E7;
    16'd40440: out <= 16'h007F;    16'd40441: out <= 16'h026E;    16'd40442: out <= 16'hF9F5;    16'd40443: out <= 16'h01F7;
    16'd40444: out <= 16'hFF04;    16'd40445: out <= 16'h0296;    16'd40446: out <= 16'h01DD;    16'd40447: out <= 16'hFFCC;
    16'd40448: out <= 16'hFE30;    16'd40449: out <= 16'h000A;    16'd40450: out <= 16'hFB1F;    16'd40451: out <= 16'h02C6;
    16'd40452: out <= 16'hFA64;    16'd40453: out <= 16'h019B;    16'd40454: out <= 16'h0125;    16'd40455: out <= 16'hFD9D;
    16'd40456: out <= 16'h0348;    16'd40457: out <= 16'h04C8;    16'd40458: out <= 16'hFA45;    16'd40459: out <= 16'h0035;
    16'd40460: out <= 16'h026B;    16'd40461: out <= 16'hFB06;    16'd40462: out <= 16'h04B8;    16'd40463: out <= 16'hFCA5;
    16'd40464: out <= 16'hF627;    16'd40465: out <= 16'h0066;    16'd40466: out <= 16'h01D6;    16'd40467: out <= 16'hFDE0;
    16'd40468: out <= 16'h03F0;    16'd40469: out <= 16'h022C;    16'd40470: out <= 16'hFA5A;    16'd40471: out <= 16'h0049;
    16'd40472: out <= 16'h0045;    16'd40473: out <= 16'hFF4B;    16'd40474: out <= 16'hFCFF;    16'd40475: out <= 16'hFB91;
    16'd40476: out <= 16'hFD54;    16'd40477: out <= 16'h0387;    16'd40478: out <= 16'hFF24;    16'd40479: out <= 16'h05B8;
    16'd40480: out <= 16'h004C;    16'd40481: out <= 16'h08F2;    16'd40482: out <= 16'hFE5F;    16'd40483: out <= 16'h07FD;
    16'd40484: out <= 16'h0647;    16'd40485: out <= 16'h0740;    16'd40486: out <= 16'h0294;    16'd40487: out <= 16'h0724;
    16'd40488: out <= 16'h03CB;    16'd40489: out <= 16'h04D7;    16'd40490: out <= 16'hFEA6;    16'd40491: out <= 16'h032D;
    16'd40492: out <= 16'hFEE2;    16'd40493: out <= 16'h0326;    16'd40494: out <= 16'h0C69;    16'd40495: out <= 16'h061A;
    16'd40496: out <= 16'h06B4;    16'd40497: out <= 16'h07A8;    16'd40498: out <= 16'h040D;    16'd40499: out <= 16'h0321;
    16'd40500: out <= 16'h0756;    16'd40501: out <= 16'h0898;    16'd40502: out <= 16'h05C3;    16'd40503: out <= 16'h07DE;
    16'd40504: out <= 16'h04A4;    16'd40505: out <= 16'hFD13;    16'd40506: out <= 16'h0201;    16'd40507: out <= 16'h001D;
    16'd40508: out <= 16'h0A50;    16'd40509: out <= 16'h048B;    16'd40510: out <= 16'hFF33;    16'd40511: out <= 16'h0348;
    16'd40512: out <= 16'h0915;    16'd40513: out <= 16'hFEDE;    16'd40514: out <= 16'h037E;    16'd40515: out <= 16'h0281;
    16'd40516: out <= 16'h03CF;    16'd40517: out <= 16'h0225;    16'd40518: out <= 16'h058D;    16'd40519: out <= 16'h025C;
    16'd40520: out <= 16'h014C;    16'd40521: out <= 16'h0631;    16'd40522: out <= 16'hFC37;    16'd40523: out <= 16'hFE3E;
    16'd40524: out <= 16'h060F;    16'd40525: out <= 16'hFEDF;    16'd40526: out <= 16'hFFE9;    16'd40527: out <= 16'h000B;
    16'd40528: out <= 16'h0162;    16'd40529: out <= 16'h028F;    16'd40530: out <= 16'h02D3;    16'd40531: out <= 16'h0241;
    16'd40532: out <= 16'h0E01;    16'd40533: out <= 16'h009D;    16'd40534: out <= 16'h0311;    16'd40535: out <= 16'h069D;
    16'd40536: out <= 16'h0515;    16'd40537: out <= 16'hFB88;    16'd40538: out <= 16'h0A3A;    16'd40539: out <= 16'hFE2E;
    16'd40540: out <= 16'h0134;    16'd40541: out <= 16'h0CA1;    16'd40542: out <= 16'h00DE;    16'd40543: out <= 16'h0587;
    16'd40544: out <= 16'h06D1;    16'd40545: out <= 16'h03A8;    16'd40546: out <= 16'h060B;    16'd40547: out <= 16'h06DA;
    16'd40548: out <= 16'hFFC5;    16'd40549: out <= 16'h0244;    16'd40550: out <= 16'h02A8;    16'd40551: out <= 16'h0690;
    16'd40552: out <= 16'h0082;    16'd40553: out <= 16'h024D;    16'd40554: out <= 16'h059C;    16'd40555: out <= 16'h0036;
    16'd40556: out <= 16'h060B;    16'd40557: out <= 16'h047E;    16'd40558: out <= 16'h0477;    16'd40559: out <= 16'h00DE;
    16'd40560: out <= 16'h006A;    16'd40561: out <= 16'hFD41;    16'd40562: out <= 16'hFF63;    16'd40563: out <= 16'hFC42;
    16'd40564: out <= 16'h06E3;    16'd40565: out <= 16'hFF2B;    16'd40566: out <= 16'h0AC7;    16'd40567: out <= 16'h01EC;
    16'd40568: out <= 16'h0340;    16'd40569: out <= 16'h00BB;    16'd40570: out <= 16'hFFE5;    16'd40571: out <= 16'h00D1;
    16'd40572: out <= 16'h0308;    16'd40573: out <= 16'h076D;    16'd40574: out <= 16'h0115;    16'd40575: out <= 16'h05C6;
    16'd40576: out <= 16'h01AA;    16'd40577: out <= 16'h0606;    16'd40578: out <= 16'h0020;    16'd40579: out <= 16'h0732;
    16'd40580: out <= 16'h00CD;    16'd40581: out <= 16'h0118;    16'd40582: out <= 16'h05E8;    16'd40583: out <= 16'h043F;
    16'd40584: out <= 16'h07B2;    16'd40585: out <= 16'h0CD6;    16'd40586: out <= 16'hFDAB;    16'd40587: out <= 16'h030A;
    16'd40588: out <= 16'h08DF;    16'd40589: out <= 16'h02FD;    16'd40590: out <= 16'h0635;    16'd40591: out <= 16'h054B;
    16'd40592: out <= 16'h06C2;    16'd40593: out <= 16'h0450;    16'd40594: out <= 16'h01F9;    16'd40595: out <= 16'h02F2;
    16'd40596: out <= 16'h0845;    16'd40597: out <= 16'h048C;    16'd40598: out <= 16'h06EE;    16'd40599: out <= 16'h0C46;
    16'd40600: out <= 16'h045A;    16'd40601: out <= 16'h03FC;    16'd40602: out <= 16'h0430;    16'd40603: out <= 16'h02F6;
    16'd40604: out <= 16'h0552;    16'd40605: out <= 16'h0268;    16'd40606: out <= 16'h044E;    16'd40607: out <= 16'h0864;
    16'd40608: out <= 16'hFE67;    16'd40609: out <= 16'h01D5;    16'd40610: out <= 16'h0739;    16'd40611: out <= 16'hFDE2;
    16'd40612: out <= 16'h02D2;    16'd40613: out <= 16'h03D3;    16'd40614: out <= 16'hFFCE;    16'd40615: out <= 16'h0452;
    16'd40616: out <= 16'h059C;    16'd40617: out <= 16'h03A4;    16'd40618: out <= 16'h0718;    16'd40619: out <= 16'h0101;
    16'd40620: out <= 16'h0413;    16'd40621: out <= 16'h0121;    16'd40622: out <= 16'h0561;    16'd40623: out <= 16'h03C7;
    16'd40624: out <= 16'hFF51;    16'd40625: out <= 16'h02CD;    16'd40626: out <= 16'h0932;    16'd40627: out <= 16'h024F;
    16'd40628: out <= 16'h01D0;    16'd40629: out <= 16'h082F;    16'd40630: out <= 16'h0421;    16'd40631: out <= 16'h040B;
    16'd40632: out <= 16'h0B38;    16'd40633: out <= 16'h02FC;    16'd40634: out <= 16'h02C1;    16'd40635: out <= 16'h03D4;
    16'd40636: out <= 16'h0193;    16'd40637: out <= 16'h07E7;    16'd40638: out <= 16'hFE6D;    16'd40639: out <= 16'h041D;
    16'd40640: out <= 16'h08E3;    16'd40641: out <= 16'h032F;    16'd40642: out <= 16'hFAF9;    16'd40643: out <= 16'h0234;
    16'd40644: out <= 16'h041F;    16'd40645: out <= 16'hFF8D;    16'd40646: out <= 16'h05B5;    16'd40647: out <= 16'h086C;
    16'd40648: out <= 16'h09AA;    16'd40649: out <= 16'h04D3;    16'd40650: out <= 16'h0637;    16'd40651: out <= 16'hFB62;
    16'd40652: out <= 16'h0957;    16'd40653: out <= 16'h03C9;    16'd40654: out <= 16'h06C8;    16'd40655: out <= 16'h0376;
    16'd40656: out <= 16'h03C2;    16'd40657: out <= 16'h08A3;    16'd40658: out <= 16'h0365;    16'd40659: out <= 16'hFE70;
    16'd40660: out <= 16'h0590;    16'd40661: out <= 16'h075F;    16'd40662: out <= 16'h036F;    16'd40663: out <= 16'h09C1;
    16'd40664: out <= 16'h05E8;    16'd40665: out <= 16'h019A;    16'd40666: out <= 16'h08B0;    16'd40667: out <= 16'h0267;
    16'd40668: out <= 16'h0A77;    16'd40669: out <= 16'h0566;    16'd40670: out <= 16'h0274;    16'd40671: out <= 16'h0775;
    16'd40672: out <= 16'h06CA;    16'd40673: out <= 16'h06D9;    16'd40674: out <= 16'h01C1;    16'd40675: out <= 16'h01C5;
    16'd40676: out <= 16'hFC4F;    16'd40677: out <= 16'hFF6F;    16'd40678: out <= 16'hFE5A;    16'd40679: out <= 16'hFF2E;
    16'd40680: out <= 16'h01E9;    16'd40681: out <= 16'h0563;    16'd40682: out <= 16'h0220;    16'd40683: out <= 16'hFEFD;
    16'd40684: out <= 16'hFECC;    16'd40685: out <= 16'h0308;    16'd40686: out <= 16'hFBFA;    16'd40687: out <= 16'h0079;
    16'd40688: out <= 16'h02ED;    16'd40689: out <= 16'h0259;    16'd40690: out <= 16'hFAD8;    16'd40691: out <= 16'h00DA;
    16'd40692: out <= 16'h00D9;    16'd40693: out <= 16'h05AF;    16'd40694: out <= 16'h0266;    16'd40695: out <= 16'h00ED;
    16'd40696: out <= 16'h0475;    16'd40697: out <= 16'h0056;    16'd40698: out <= 16'h02AB;    16'd40699: out <= 16'h0034;
    16'd40700: out <= 16'hFECB;    16'd40701: out <= 16'hFF02;    16'd40702: out <= 16'hFF49;    16'd40703: out <= 16'hF959;
    16'd40704: out <= 16'h00A4;    16'd40705: out <= 16'h021E;    16'd40706: out <= 16'h01F6;    16'd40707: out <= 16'h05E6;
    16'd40708: out <= 16'hFEA5;    16'd40709: out <= 16'h0311;    16'd40710: out <= 16'h01E4;    16'd40711: out <= 16'h0155;
    16'd40712: out <= 16'hFBE3;    16'd40713: out <= 16'h04AD;    16'd40714: out <= 16'hFE6F;    16'd40715: out <= 16'h0302;
    16'd40716: out <= 16'hF840;    16'd40717: out <= 16'h0610;    16'd40718: out <= 16'hF797;    16'd40719: out <= 16'h0490;
    16'd40720: out <= 16'hFC0C;    16'd40721: out <= 16'hFA84;    16'd40722: out <= 16'hF977;    16'd40723: out <= 16'hFD24;
    16'd40724: out <= 16'hFD59;    16'd40725: out <= 16'hF951;    16'd40726: out <= 16'hFFC4;    16'd40727: out <= 16'h0248;
    16'd40728: out <= 16'h0343;    16'd40729: out <= 16'h00C0;    16'd40730: out <= 16'h059C;    16'd40731: out <= 16'h0220;
    16'd40732: out <= 16'h0061;    16'd40733: out <= 16'hFBD4;    16'd40734: out <= 16'h0190;    16'd40735: out <= 16'h03D1;
    16'd40736: out <= 16'h0B31;    16'd40737: out <= 16'hFBE9;    16'd40738: out <= 16'hFC02;    16'd40739: out <= 16'h0AC0;
    16'd40740: out <= 16'h039A;    16'd40741: out <= 16'hFFB7;    16'd40742: out <= 16'h1091;    16'd40743: out <= 16'hFF62;
    16'd40744: out <= 16'hFB3C;    16'd40745: out <= 16'hFFD7;    16'd40746: out <= 16'h040B;    16'd40747: out <= 16'hFAFB;
    16'd40748: out <= 16'h03A0;    16'd40749: out <= 16'h0372;    16'd40750: out <= 16'h03D1;    16'd40751: out <= 16'h0517;
    16'd40752: out <= 16'h02A2;    16'd40753: out <= 16'hFEEA;    16'd40754: out <= 16'h0474;    16'd40755: out <= 16'hFF5E;
    16'd40756: out <= 16'h031B;    16'd40757: out <= 16'hFFFC;    16'd40758: out <= 16'h043A;    16'd40759: out <= 16'h0551;
    16'd40760: out <= 16'h01C7;    16'd40761: out <= 16'h05BF;    16'd40762: out <= 16'h001D;    16'd40763: out <= 16'h020D;
    16'd40764: out <= 16'h039E;    16'd40765: out <= 16'h04A5;    16'd40766: out <= 16'h083C;    16'd40767: out <= 16'h016A;
    16'd40768: out <= 16'hFA8F;    16'd40769: out <= 16'h0708;    16'd40770: out <= 16'h020A;    16'd40771: out <= 16'h012F;
    16'd40772: out <= 16'h0416;    16'd40773: out <= 16'h01BC;    16'd40774: out <= 16'h083F;    16'd40775: out <= 16'h0470;
    16'd40776: out <= 16'hFEDE;    16'd40777: out <= 16'hFB57;    16'd40778: out <= 16'h09CF;    16'd40779: out <= 16'hFA70;
    16'd40780: out <= 16'h0865;    16'd40781: out <= 16'h0726;    16'd40782: out <= 16'h0314;    16'd40783: out <= 16'h01AA;
    16'd40784: out <= 16'h04DD;    16'd40785: out <= 16'h063D;    16'd40786: out <= 16'h08B4;    16'd40787: out <= 16'hFA7C;
    16'd40788: out <= 16'h0485;    16'd40789: out <= 16'h0749;    16'd40790: out <= 16'h05C0;    16'd40791: out <= 16'h00CA;
    16'd40792: out <= 16'h02F3;    16'd40793: out <= 16'h03CC;    16'd40794: out <= 16'hFEF5;    16'd40795: out <= 16'hF8C3;
    16'd40796: out <= 16'h03E3;    16'd40797: out <= 16'h08A0;    16'd40798: out <= 16'h06EE;    16'd40799: out <= 16'h052D;
    16'd40800: out <= 16'h0125;    16'd40801: out <= 16'h0250;    16'd40802: out <= 16'h013A;    16'd40803: out <= 16'h079E;
    16'd40804: out <= 16'h0163;    16'd40805: out <= 16'h0337;    16'd40806: out <= 16'h00A1;    16'd40807: out <= 16'h03E9;
    16'd40808: out <= 16'h0413;    16'd40809: out <= 16'h05E3;    16'd40810: out <= 16'h09D0;    16'd40811: out <= 16'h01B2;
    16'd40812: out <= 16'h0A29;    16'd40813: out <= 16'h07E9;    16'd40814: out <= 16'hFCB4;    16'd40815: out <= 16'hFBA1;
    16'd40816: out <= 16'h00CE;    16'd40817: out <= 16'h087C;    16'd40818: out <= 16'h042E;    16'd40819: out <= 16'h036A;
    16'd40820: out <= 16'h0877;    16'd40821: out <= 16'h0265;    16'd40822: out <= 16'hFAC9;    16'd40823: out <= 16'h05FD;
    16'd40824: out <= 16'h00EB;    16'd40825: out <= 16'h0620;    16'd40826: out <= 16'h02F7;    16'd40827: out <= 16'h074C;
    16'd40828: out <= 16'h0119;    16'd40829: out <= 16'h020C;    16'd40830: out <= 16'h055B;    16'd40831: out <= 16'hFFC8;
    16'd40832: out <= 16'hFF40;    16'd40833: out <= 16'h03D2;    16'd40834: out <= 16'h051F;    16'd40835: out <= 16'h00DA;
    16'd40836: out <= 16'h0478;    16'd40837: out <= 16'h0311;    16'd40838: out <= 16'h01DD;    16'd40839: out <= 16'h0890;
    16'd40840: out <= 16'h05AE;    16'd40841: out <= 16'h0103;    16'd40842: out <= 16'h05BD;    16'd40843: out <= 16'hFCB3;
    16'd40844: out <= 16'h0805;    16'd40845: out <= 16'h069C;    16'd40846: out <= 16'h0719;    16'd40847: out <= 16'h0112;
    16'd40848: out <= 16'h046F;    16'd40849: out <= 16'h06F3;    16'd40850: out <= 16'h0667;    16'd40851: out <= 16'h01AA;
    16'd40852: out <= 16'hFF9A;    16'd40853: out <= 16'h059F;    16'd40854: out <= 16'h0332;    16'd40855: out <= 16'h064F;
    16'd40856: out <= 16'h034B;    16'd40857: out <= 16'h04F0;    16'd40858: out <= 16'hFD20;    16'd40859: out <= 16'h0A59;
    16'd40860: out <= 16'h0616;    16'd40861: out <= 16'h0369;    16'd40862: out <= 16'h04C8;    16'd40863: out <= 16'h0067;
    16'd40864: out <= 16'h070E;    16'd40865: out <= 16'h078F;    16'd40866: out <= 16'h015D;    16'd40867: out <= 16'hFF64;
    16'd40868: out <= 16'h0219;    16'd40869: out <= 16'h0455;    16'd40870: out <= 16'h0077;    16'd40871: out <= 16'h064B;
    16'd40872: out <= 16'hFD46;    16'd40873: out <= 16'hFFB1;    16'd40874: out <= 16'h0544;    16'd40875: out <= 16'h022B;
    16'd40876: out <= 16'h01A5;    16'd40877: out <= 16'h05E0;    16'd40878: out <= 16'h0711;    16'd40879: out <= 16'h06C2;
    16'd40880: out <= 16'h0549;    16'd40881: out <= 16'h081A;    16'd40882: out <= 16'h06FD;    16'd40883: out <= 16'h037B;
    16'd40884: out <= 16'hFD2E;    16'd40885: out <= 16'h0333;    16'd40886: out <= 16'h01F2;    16'd40887: out <= 16'h043E;
    16'd40888: out <= 16'h014E;    16'd40889: out <= 16'hFE92;    16'd40890: out <= 16'h00D9;    16'd40891: out <= 16'h02F3;
    16'd40892: out <= 16'h0668;    16'd40893: out <= 16'h0277;    16'd40894: out <= 16'h0831;    16'd40895: out <= 16'h08C5;
    16'd40896: out <= 16'h071F;    16'd40897: out <= 16'h0292;    16'd40898: out <= 16'h021D;    16'd40899: out <= 16'h0054;
    16'd40900: out <= 16'h048F;    16'd40901: out <= 16'h0507;    16'd40902: out <= 16'hFF8F;    16'd40903: out <= 16'h009E;
    16'd40904: out <= 16'h0AC0;    16'd40905: out <= 16'h0608;    16'd40906: out <= 16'h009E;    16'd40907: out <= 16'hFDFE;
    16'd40908: out <= 16'hFB9B;    16'd40909: out <= 16'h0A6C;    16'd40910: out <= 16'h00AC;    16'd40911: out <= 16'h00EE;
    16'd40912: out <= 16'h057B;    16'd40913: out <= 16'h056E;    16'd40914: out <= 16'h019E;    16'd40915: out <= 16'h059B;
    16'd40916: out <= 16'h0805;    16'd40917: out <= 16'h00A5;    16'd40918: out <= 16'h050F;    16'd40919: out <= 16'h09F1;
    16'd40920: out <= 16'hFECF;    16'd40921: out <= 16'h05E8;    16'd40922: out <= 16'hFF69;    16'd40923: out <= 16'h0083;
    16'd40924: out <= 16'h0400;    16'd40925: out <= 16'hFD8D;    16'd40926: out <= 16'h03D8;    16'd40927: out <= 16'h03D2;
    16'd40928: out <= 16'h0284;    16'd40929: out <= 16'hFA46;    16'd40930: out <= 16'h04D9;    16'd40931: out <= 16'hFED5;
    16'd40932: out <= 16'hFAB6;    16'd40933: out <= 16'hFC6C;    16'd40934: out <= 16'hF795;    16'd40935: out <= 16'hF8B0;
    16'd40936: out <= 16'h017E;    16'd40937: out <= 16'h03D2;    16'd40938: out <= 16'h004E;    16'd40939: out <= 16'h0088;
    16'd40940: out <= 16'hF7DD;    16'd40941: out <= 16'hFB8B;    16'd40942: out <= 16'h039C;    16'd40943: out <= 16'hFBEC;
    16'd40944: out <= 16'h00F9;    16'd40945: out <= 16'h000A;    16'd40946: out <= 16'h01DB;    16'd40947: out <= 16'h0166;
    16'd40948: out <= 16'h07F0;    16'd40949: out <= 16'hFC10;    16'd40950: out <= 16'hFD6C;    16'd40951: out <= 16'hFE84;
    16'd40952: out <= 16'hF757;    16'd40953: out <= 16'h00B2;    16'd40954: out <= 16'h0295;    16'd40955: out <= 16'h00DE;
    16'd40956: out <= 16'hFE45;    16'd40957: out <= 16'hFC14;    16'd40958: out <= 16'hFDE7;    16'd40959: out <= 16'h0629;
    16'd40960: out <= 16'hFDD7;    16'd40961: out <= 16'h03CC;    16'd40962: out <= 16'hFC20;    16'd40963: out <= 16'hFE6E;
    16'd40964: out <= 16'h04B7;    16'd40965: out <= 16'hFC55;    16'd40966: out <= 16'h031E;    16'd40967: out <= 16'h02B0;
    16'd40968: out <= 16'h0769;    16'd40969: out <= 16'h01D0;    16'd40970: out <= 16'h082C;    16'd40971: out <= 16'h064B;
    16'd40972: out <= 16'hFE2B;    16'd40973: out <= 16'h04FB;    16'd40974: out <= 16'hFD16;    16'd40975: out <= 16'h0472;
    16'd40976: out <= 16'h0248;    16'd40977: out <= 16'hFFF1;    16'd40978: out <= 16'h0372;    16'd40979: out <= 16'h0352;
    16'd40980: out <= 16'h0950;    16'd40981: out <= 16'h00A0;    16'd40982: out <= 16'h024D;    16'd40983: out <= 16'hFFFD;
    16'd40984: out <= 16'h021C;    16'd40985: out <= 16'h096D;    16'd40986: out <= 16'h0045;    16'd40987: out <= 16'hFD5F;
    16'd40988: out <= 16'h01FE;    16'd40989: out <= 16'hFB90;    16'd40990: out <= 16'h0377;    16'd40991: out <= 16'h01A3;
    16'd40992: out <= 16'h079F;    16'd40993: out <= 16'hFFF2;    16'd40994: out <= 16'h0445;    16'd40995: out <= 16'h03BD;
    16'd40996: out <= 16'h01E0;    16'd40997: out <= 16'hFF1E;    16'd40998: out <= 16'hFE81;    16'd40999: out <= 16'h05D1;
    16'd41000: out <= 16'h0BBB;    16'd41001: out <= 16'h0383;    16'd41002: out <= 16'h05B0;    16'd41003: out <= 16'h06B5;
    16'd41004: out <= 16'h02E8;    16'd41005: out <= 16'h03DA;    16'd41006: out <= 16'h0016;    16'd41007: out <= 16'h0346;
    16'd41008: out <= 16'h0456;    16'd41009: out <= 16'h04E6;    16'd41010: out <= 16'hFBD6;    16'd41011: out <= 16'hFC82;
    16'd41012: out <= 16'hFDB4;    16'd41013: out <= 16'h083C;    16'd41014: out <= 16'h0C07;    16'd41015: out <= 16'hFF55;
    16'd41016: out <= 16'h069E;    16'd41017: out <= 16'h03C5;    16'd41018: out <= 16'h0B32;    16'd41019: out <= 16'h08E0;
    16'd41020: out <= 16'h01E8;    16'd41021: out <= 16'h00BD;    16'd41022: out <= 16'h0548;    16'd41023: out <= 16'hFFC5;
    16'd41024: out <= 16'h0253;    16'd41025: out <= 16'h09F8;    16'd41026: out <= 16'h05D9;    16'd41027: out <= 16'hFB78;
    16'd41028: out <= 16'h0407;    16'd41029: out <= 16'h0222;    16'd41030: out <= 16'h0046;    16'd41031: out <= 16'h0570;
    16'd41032: out <= 16'h01A9;    16'd41033: out <= 16'h0884;    16'd41034: out <= 16'h03DE;    16'd41035: out <= 16'h0AE8;
    16'd41036: out <= 16'h04B5;    16'd41037: out <= 16'h0097;    16'd41038: out <= 16'h002B;    16'd41039: out <= 16'h03C5;
    16'd41040: out <= 16'hFF4D;    16'd41041: out <= 16'h0408;    16'd41042: out <= 16'h073B;    16'd41043: out <= 16'hFA85;
    16'd41044: out <= 16'h07B4;    16'd41045: out <= 16'h0343;    16'd41046: out <= 16'h058A;    16'd41047: out <= 16'hFD5C;
    16'd41048: out <= 16'h0212;    16'd41049: out <= 16'hFC9C;    16'd41050: out <= 16'h057D;    16'd41051: out <= 16'h040E;
    16'd41052: out <= 16'h0186;    16'd41053: out <= 16'h03D5;    16'd41054: out <= 16'hFECD;    16'd41055: out <= 16'h0722;
    16'd41056: out <= 16'h0773;    16'd41057: out <= 16'h0A02;    16'd41058: out <= 16'h08EC;    16'd41059: out <= 16'h02A7;
    16'd41060: out <= 16'h03EE;    16'd41061: out <= 16'h0384;    16'd41062: out <= 16'h0886;    16'd41063: out <= 16'hFF68;
    16'd41064: out <= 16'h0153;    16'd41065: out <= 16'h0A91;    16'd41066: out <= 16'h06D6;    16'd41067: out <= 16'h0849;
    16'd41068: out <= 16'hF8E9;    16'd41069: out <= 16'hFE72;    16'd41070: out <= 16'h0048;    16'd41071: out <= 16'hFEB4;
    16'd41072: out <= 16'hFED5;    16'd41073: out <= 16'hFE9A;    16'd41074: out <= 16'h0449;    16'd41075: out <= 16'hFFE4;
    16'd41076: out <= 16'h05D5;    16'd41077: out <= 16'h0477;    16'd41078: out <= 16'h03AB;    16'd41079: out <= 16'h0644;
    16'd41080: out <= 16'h0511;    16'd41081: out <= 16'h01E9;    16'd41082: out <= 16'h037F;    16'd41083: out <= 16'h0214;
    16'd41084: out <= 16'h0A35;    16'd41085: out <= 16'hFF83;    16'd41086: out <= 16'h023A;    16'd41087: out <= 16'h0D76;
    16'd41088: out <= 16'h07A0;    16'd41089: out <= 16'h0792;    16'd41090: out <= 16'h03EC;    16'd41091: out <= 16'h00D6;
    16'd41092: out <= 16'h01F5;    16'd41093: out <= 16'h017D;    16'd41094: out <= 16'h0198;    16'd41095: out <= 16'h083C;
    16'd41096: out <= 16'hFB0C;    16'd41097: out <= 16'h051A;    16'd41098: out <= 16'h05A4;    16'd41099: out <= 16'hFEB8;
    16'd41100: out <= 16'h001E;    16'd41101: out <= 16'h076D;    16'd41102: out <= 16'h068B;    16'd41103: out <= 16'h01EC;
    16'd41104: out <= 16'h05A9;    16'd41105: out <= 16'h0786;    16'd41106: out <= 16'h004D;    16'd41107: out <= 16'hFF0C;
    16'd41108: out <= 16'h0806;    16'd41109: out <= 16'h02BC;    16'd41110: out <= 16'h09C4;    16'd41111: out <= 16'h07B0;
    16'd41112: out <= 16'h03F5;    16'd41113: out <= 16'h0290;    16'd41114: out <= 16'h0737;    16'd41115: out <= 16'h0408;
    16'd41116: out <= 16'hFCED;    16'd41117: out <= 16'hFFA2;    16'd41118: out <= 16'h0256;    16'd41119: out <= 16'h035F;
    16'd41120: out <= 16'h0290;    16'd41121: out <= 16'h0938;    16'd41122: out <= 16'h0012;    16'd41123: out <= 16'h0809;
    16'd41124: out <= 16'h045F;    16'd41125: out <= 16'h096B;    16'd41126: out <= 16'h0046;    16'd41127: out <= 16'h0579;
    16'd41128: out <= 16'h06AB;    16'd41129: out <= 16'h03A8;    16'd41130: out <= 16'h0349;    16'd41131: out <= 16'h07B1;
    16'd41132: out <= 16'h077D;    16'd41133: out <= 16'h0228;    16'd41134: out <= 16'h0232;    16'd41135: out <= 16'h057E;
    16'd41136: out <= 16'h0466;    16'd41137: out <= 16'h0621;    16'd41138: out <= 16'h02C8;    16'd41139: out <= 16'h04B5;
    16'd41140: out <= 16'h00F4;    16'd41141: out <= 16'h0632;    16'd41142: out <= 16'h0324;    16'd41143: out <= 16'h0255;
    16'd41144: out <= 16'h0A57;    16'd41145: out <= 16'h07F0;    16'd41146: out <= 16'h0771;    16'd41147: out <= 16'h059D;
    16'd41148: out <= 16'h07DE;    16'd41149: out <= 16'h00B4;    16'd41150: out <= 16'h0AB5;    16'd41151: out <= 16'h02BE;
    16'd41152: out <= 16'h04D6;    16'd41153: out <= 16'h09B9;    16'd41154: out <= 16'h0779;    16'd41155: out <= 16'h07A8;
    16'd41156: out <= 16'h05C1;    16'd41157: out <= 16'hFEE9;    16'd41158: out <= 16'h0496;    16'd41159: out <= 16'h0349;
    16'd41160: out <= 16'h014C;    16'd41161: out <= 16'h0590;    16'd41162: out <= 16'h062E;    16'd41163: out <= 16'h0B1E;
    16'd41164: out <= 16'h04F6;    16'd41165: out <= 16'h08EC;    16'd41166: out <= 16'hFD01;    16'd41167: out <= 16'h03E8;
    16'd41168: out <= 16'h02C5;    16'd41169: out <= 16'h01A1;    16'd41170: out <= 16'hFF4F;    16'd41171: out <= 16'h04CA;
    16'd41172: out <= 16'h03D2;    16'd41173: out <= 16'hFC1E;    16'd41174: out <= 16'hFFDC;    16'd41175: out <= 16'h0289;
    16'd41176: out <= 16'h04F1;    16'd41177: out <= 16'h021A;    16'd41178: out <= 16'h05DD;    16'd41179: out <= 16'h03DD;
    16'd41180: out <= 16'h07C7;    16'd41181: out <= 16'h04B0;    16'd41182: out <= 16'h056C;    16'd41183: out <= 16'h01A2;
    16'd41184: out <= 16'hFDAE;    16'd41185: out <= 16'h0954;    16'd41186: out <= 16'h0944;    16'd41187: out <= 16'h04B5;
    16'd41188: out <= 16'hFC2A;    16'd41189: out <= 16'hFFC2;    16'd41190: out <= 16'h0819;    16'd41191: out <= 16'hFAC2;
    16'd41192: out <= 16'hFB41;    16'd41193: out <= 16'hFEAE;    16'd41194: out <= 16'hFEF5;    16'd41195: out <= 16'hFBA7;
    16'd41196: out <= 16'hFF05;    16'd41197: out <= 16'h0186;    16'd41198: out <= 16'h0247;    16'd41199: out <= 16'hFC32;
    16'd41200: out <= 16'hFFFB;    16'd41201: out <= 16'hFC7A;    16'd41202: out <= 16'h0ACC;    16'd41203: out <= 16'h0383;
    16'd41204: out <= 16'hFF78;    16'd41205: out <= 16'h02BF;    16'd41206: out <= 16'h07E6;    16'd41207: out <= 16'h0141;
    16'd41208: out <= 16'hFAB9;    16'd41209: out <= 16'hFC8D;    16'd41210: out <= 16'h038D;    16'd41211: out <= 16'hFD0A;
    16'd41212: out <= 16'h00CB;    16'd41213: out <= 16'h0617;    16'd41214: out <= 16'hFA9E;    16'd41215: out <= 16'hFF09;
    16'd41216: out <= 16'hFF1C;    16'd41217: out <= 16'h0256;    16'd41218: out <= 16'h014A;    16'd41219: out <= 16'hFBAB;
    16'd41220: out <= 16'h05A0;    16'd41221: out <= 16'h0102;    16'd41222: out <= 16'hFC92;    16'd41223: out <= 16'h0697;
    16'd41224: out <= 16'h034C;    16'd41225: out <= 16'hFD17;    16'd41226: out <= 16'hFF83;    16'd41227: out <= 16'h0559;
    16'd41228: out <= 16'h0007;    16'd41229: out <= 16'hFF87;    16'd41230: out <= 16'h0349;    16'd41231: out <= 16'h00BC;
    16'd41232: out <= 16'h0485;    16'd41233: out <= 16'h0406;    16'd41234: out <= 16'h0460;    16'd41235: out <= 16'h07B5;
    16'd41236: out <= 16'h011E;    16'd41237: out <= 16'hFD79;    16'd41238: out <= 16'h001F;    16'd41239: out <= 16'hFDBF;
    16'd41240: out <= 16'hF9C2;    16'd41241: out <= 16'h0001;    16'd41242: out <= 16'hFE38;    16'd41243: out <= 16'h08C8;
    16'd41244: out <= 16'h0119;    16'd41245: out <= 16'h01C0;    16'd41246: out <= 16'h03B9;    16'd41247: out <= 16'h0173;
    16'd41248: out <= 16'h09D3;    16'd41249: out <= 16'hFE47;    16'd41250: out <= 16'hFFCB;    16'd41251: out <= 16'h0391;
    16'd41252: out <= 16'h0533;    16'd41253: out <= 16'h0BBE;    16'd41254: out <= 16'h0371;    16'd41255: out <= 16'h08F2;
    16'd41256: out <= 16'h03B9;    16'd41257: out <= 16'h03DB;    16'd41258: out <= 16'h04CB;    16'd41259: out <= 16'hFDF1;
    16'd41260: out <= 16'h01FA;    16'd41261: out <= 16'h031E;    16'd41262: out <= 16'h058B;    16'd41263: out <= 16'hFE30;
    16'd41264: out <= 16'h00B2;    16'd41265: out <= 16'h0205;    16'd41266: out <= 16'h05EF;    16'd41267: out <= 16'h004A;
    16'd41268: out <= 16'hFE9F;    16'd41269: out <= 16'hFD2B;    16'd41270: out <= 16'hFD9C;    16'd41271: out <= 16'h08E2;
    16'd41272: out <= 16'h05B3;    16'd41273: out <= 16'h02F0;    16'd41274: out <= 16'h07F1;    16'd41275: out <= 16'h0258;
    16'd41276: out <= 16'hFDA2;    16'd41277: out <= 16'h0277;    16'd41278: out <= 16'h0060;    16'd41279: out <= 16'hFEAB;
    16'd41280: out <= 16'hFD61;    16'd41281: out <= 16'h04E3;    16'd41282: out <= 16'h0640;    16'd41283: out <= 16'hFE9E;
    16'd41284: out <= 16'hFF29;    16'd41285: out <= 16'h0311;    16'd41286: out <= 16'h0428;    16'd41287: out <= 16'h0266;
    16'd41288: out <= 16'h00AA;    16'd41289: out <= 16'hFDCE;    16'd41290: out <= 16'h02BE;    16'd41291: out <= 16'h001A;
    16'd41292: out <= 16'h05E1;    16'd41293: out <= 16'h03C9;    16'd41294: out <= 16'h0392;    16'd41295: out <= 16'h03B8;
    16'd41296: out <= 16'h000E;    16'd41297: out <= 16'h0292;    16'd41298: out <= 16'hFEDA;    16'd41299: out <= 16'h0288;
    16'd41300: out <= 16'h036C;    16'd41301: out <= 16'h090B;    16'd41302: out <= 16'hFF8C;    16'd41303: out <= 16'hFE1D;
    16'd41304: out <= 16'h02AB;    16'd41305: out <= 16'h0921;    16'd41306: out <= 16'h01C8;    16'd41307: out <= 16'h0229;
    16'd41308: out <= 16'hFF53;    16'd41309: out <= 16'hFDA8;    16'd41310: out <= 16'h034B;    16'd41311: out <= 16'h047C;
    16'd41312: out <= 16'h056B;    16'd41313: out <= 16'h03DF;    16'd41314: out <= 16'h09BE;    16'd41315: out <= 16'h09E2;
    16'd41316: out <= 16'h072C;    16'd41317: out <= 16'h00C6;    16'd41318: out <= 16'h062E;    16'd41319: out <= 16'h020B;
    16'd41320: out <= 16'h088B;    16'd41321: out <= 16'h0634;    16'd41322: out <= 16'h03F0;    16'd41323: out <= 16'h01B5;
    16'd41324: out <= 16'h03EF;    16'd41325: out <= 16'h0345;    16'd41326: out <= 16'h02EC;    16'd41327: out <= 16'h06C0;
    16'd41328: out <= 16'h0825;    16'd41329: out <= 16'h00F3;    16'd41330: out <= 16'h0443;    16'd41331: out <= 16'h0307;
    16'd41332: out <= 16'h0127;    16'd41333: out <= 16'h060F;    16'd41334: out <= 16'h070C;    16'd41335: out <= 16'h0814;
    16'd41336: out <= 16'h0A35;    16'd41337: out <= 16'h0973;    16'd41338: out <= 16'h015A;    16'd41339: out <= 16'h00C7;
    16'd41340: out <= 16'h02A8;    16'd41341: out <= 16'h0377;    16'd41342: out <= 16'h01DE;    16'd41343: out <= 16'h099F;
    16'd41344: out <= 16'h045D;    16'd41345: out <= 16'h04CD;    16'd41346: out <= 16'h0224;    16'd41347: out <= 16'h0B4C;
    16'd41348: out <= 16'hFF04;    16'd41349: out <= 16'h096A;    16'd41350: out <= 16'h02AC;    16'd41351: out <= 16'h0C1F;
    16'd41352: out <= 16'h02B8;    16'd41353: out <= 16'h05D9;    16'd41354: out <= 16'h032F;    16'd41355: out <= 16'h0459;
    16'd41356: out <= 16'hFEC4;    16'd41357: out <= 16'h04D0;    16'd41358: out <= 16'h023F;    16'd41359: out <= 16'h04C2;
    16'd41360: out <= 16'h08CB;    16'd41361: out <= 16'h0353;    16'd41362: out <= 16'h0F5D;    16'd41363: out <= 16'h08A6;
    16'd41364: out <= 16'hFC05;    16'd41365: out <= 16'h0496;    16'd41366: out <= 16'h01EE;    16'd41367: out <= 16'h070C;
    16'd41368: out <= 16'h0644;    16'd41369: out <= 16'h080D;    16'd41370: out <= 16'h003F;    16'd41371: out <= 16'h065C;
    16'd41372: out <= 16'hFFBE;    16'd41373: out <= 16'h0AEA;    16'd41374: out <= 16'h06FD;    16'd41375: out <= 16'h0A53;
    16'd41376: out <= 16'hFB4B;    16'd41377: out <= 16'hFDF3;    16'd41378: out <= 16'h066A;    16'd41379: out <= 16'h0497;
    16'd41380: out <= 16'h001E;    16'd41381: out <= 16'h0CFD;    16'd41382: out <= 16'hFEC5;    16'd41383: out <= 16'h0504;
    16'd41384: out <= 16'h00EC;    16'd41385: out <= 16'hFDDB;    16'd41386: out <= 16'h004F;    16'd41387: out <= 16'h0802;
    16'd41388: out <= 16'h004D;    16'd41389: out <= 16'h04D3;    16'd41390: out <= 16'h0892;    16'd41391: out <= 16'hFFEA;
    16'd41392: out <= 16'hFE08;    16'd41393: out <= 16'h051B;    16'd41394: out <= 16'h0409;    16'd41395: out <= 16'hFBBC;
    16'd41396: out <= 16'h0710;    16'd41397: out <= 16'h0359;    16'd41398: out <= 16'h037B;    16'd41399: out <= 16'h05C9;
    16'd41400: out <= 16'h032B;    16'd41401: out <= 16'h04B6;    16'd41402: out <= 16'h0899;    16'd41403: out <= 16'h0254;
    16'd41404: out <= 16'hFE44;    16'd41405: out <= 16'hFA3C;    16'd41406: out <= 16'h017C;    16'd41407: out <= 16'h0488;
    16'd41408: out <= 16'h0297;    16'd41409: out <= 16'h055E;    16'd41410: out <= 16'h08D4;    16'd41411: out <= 16'hFB6E;
    16'd41412: out <= 16'h01CD;    16'd41413: out <= 16'h0646;    16'd41414: out <= 16'h00E9;    16'd41415: out <= 16'hFF24;
    16'd41416: out <= 16'h02DE;    16'd41417: out <= 16'h00F1;    16'd41418: out <= 16'h0140;    16'd41419: out <= 16'h037B;
    16'd41420: out <= 16'h06B2;    16'd41421: out <= 16'h03DE;    16'd41422: out <= 16'h089F;    16'd41423: out <= 16'h02B2;
    16'd41424: out <= 16'h041E;    16'd41425: out <= 16'h052C;    16'd41426: out <= 16'h00E7;    16'd41427: out <= 16'h03C2;
    16'd41428: out <= 16'h086A;    16'd41429: out <= 16'h00E8;    16'd41430: out <= 16'h0527;    16'd41431: out <= 16'h0168;
    16'd41432: out <= 16'hFC69;    16'd41433: out <= 16'h05DF;    16'd41434: out <= 16'h0549;    16'd41435: out <= 16'h0656;
    16'd41436: out <= 16'h00A4;    16'd41437: out <= 16'h0537;    16'd41438: out <= 16'h00E8;    16'd41439: out <= 16'h02D9;
    16'd41440: out <= 16'h06F9;    16'd41441: out <= 16'hFE47;    16'd41442: out <= 16'hFE5C;    16'd41443: out <= 16'h0054;
    16'd41444: out <= 16'h00A4;    16'd41445: out <= 16'hFE5A;    16'd41446: out <= 16'hFF85;    16'd41447: out <= 16'h0461;
    16'd41448: out <= 16'hFE13;    16'd41449: out <= 16'hFF13;    16'd41450: out <= 16'hF952;    16'd41451: out <= 16'hFE8D;
    16'd41452: out <= 16'h01B7;    16'd41453: out <= 16'hFDCE;    16'd41454: out <= 16'h024B;    16'd41455: out <= 16'hFD0D;
    16'd41456: out <= 16'hFD79;    16'd41457: out <= 16'hFF52;    16'd41458: out <= 16'h06A2;    16'd41459: out <= 16'hFCF6;
    16'd41460: out <= 16'h059C;    16'd41461: out <= 16'h01F0;    16'd41462: out <= 16'h0545;    16'd41463: out <= 16'h017F;
    16'd41464: out <= 16'hFB32;    16'd41465: out <= 16'hFC27;    16'd41466: out <= 16'h05D3;    16'd41467: out <= 16'h064E;
    16'd41468: out <= 16'hFFC5;    16'd41469: out <= 16'h0035;    16'd41470: out <= 16'h0125;    16'd41471: out <= 16'hFF36;
    16'd41472: out <= 16'h008D;    16'd41473: out <= 16'hFF8C;    16'd41474: out <= 16'h05A1;    16'd41475: out <= 16'hFDB8;
    16'd41476: out <= 16'h0871;    16'd41477: out <= 16'h0075;    16'd41478: out <= 16'h00AE;    16'd41479: out <= 16'h0333;
    16'd41480: out <= 16'h0194;    16'd41481: out <= 16'hFD6B;    16'd41482: out <= 16'hFDD8;    16'd41483: out <= 16'hFB41;
    16'd41484: out <= 16'h0023;    16'd41485: out <= 16'h0726;    16'd41486: out <= 16'h01E3;    16'd41487: out <= 16'hFE3B;
    16'd41488: out <= 16'hFF10;    16'd41489: out <= 16'h02E4;    16'd41490: out <= 16'h059E;    16'd41491: out <= 16'h0349;
    16'd41492: out <= 16'hFFC5;    16'd41493: out <= 16'h07DB;    16'd41494: out <= 16'hFE35;    16'd41495: out <= 16'hF8F3;
    16'd41496: out <= 16'h0076;    16'd41497: out <= 16'h01F3;    16'd41498: out <= 16'h00B8;    16'd41499: out <= 16'hFE98;
    16'd41500: out <= 16'hFF20;    16'd41501: out <= 16'h0336;    16'd41502: out <= 16'h0AFF;    16'd41503: out <= 16'h0258;
    16'd41504: out <= 16'h008E;    16'd41505: out <= 16'h0725;    16'd41506: out <= 16'h0363;    16'd41507: out <= 16'h0173;
    16'd41508: out <= 16'h019A;    16'd41509: out <= 16'hFD5B;    16'd41510: out <= 16'h0047;    16'd41511: out <= 16'h0467;
    16'd41512: out <= 16'h0694;    16'd41513: out <= 16'hFD38;    16'd41514: out <= 16'h0019;    16'd41515: out <= 16'hFF34;
    16'd41516: out <= 16'h014C;    16'd41517: out <= 16'hFE3D;    16'd41518: out <= 16'h0848;    16'd41519: out <= 16'h070A;
    16'd41520: out <= 16'h0A52;    16'd41521: out <= 16'h0088;    16'd41522: out <= 16'h02E8;    16'd41523: out <= 16'h02A4;
    16'd41524: out <= 16'h0A4F;    16'd41525: out <= 16'h03B7;    16'd41526: out <= 16'h09D9;    16'd41527: out <= 16'h080F;
    16'd41528: out <= 16'h0B85;    16'd41529: out <= 16'h03E2;    16'd41530: out <= 16'h0350;    16'd41531: out <= 16'h098E;
    16'd41532: out <= 16'h0986;    16'd41533: out <= 16'hF8E2;    16'd41534: out <= 16'hFBD2;    16'd41535: out <= 16'hFE84;
    16'd41536: out <= 16'h03A8;    16'd41537: out <= 16'h064A;    16'd41538: out <= 16'hFFC1;    16'd41539: out <= 16'h031F;
    16'd41540: out <= 16'h0096;    16'd41541: out <= 16'h0156;    16'd41542: out <= 16'hFF81;    16'd41543: out <= 16'h0796;
    16'd41544: out <= 16'h0155;    16'd41545: out <= 16'hFC5A;    16'd41546: out <= 16'h02E6;    16'd41547: out <= 16'hFF59;
    16'd41548: out <= 16'h0250;    16'd41549: out <= 16'h0424;    16'd41550: out <= 16'h01FF;    16'd41551: out <= 16'h014E;
    16'd41552: out <= 16'h034F;    16'd41553: out <= 16'hFE12;    16'd41554: out <= 16'h0396;    16'd41555: out <= 16'h0321;
    16'd41556: out <= 16'hFBA3;    16'd41557: out <= 16'hF8BE;    16'd41558: out <= 16'h0A90;    16'd41559: out <= 16'h02CE;
    16'd41560: out <= 16'h06F8;    16'd41561: out <= 16'h020D;    16'd41562: out <= 16'h0138;    16'd41563: out <= 16'h022E;
    16'd41564: out <= 16'h0275;    16'd41565: out <= 16'h037E;    16'd41566: out <= 16'h0A70;    16'd41567: out <= 16'hFEC2;
    16'd41568: out <= 16'hFD06;    16'd41569: out <= 16'h0402;    16'd41570: out <= 16'hFD67;    16'd41571: out <= 16'h03B3;
    16'd41572: out <= 16'h073B;    16'd41573: out <= 16'h05BE;    16'd41574: out <= 16'h071D;    16'd41575: out <= 16'h0461;
    16'd41576: out <= 16'hFEDA;    16'd41577: out <= 16'h06C2;    16'd41578: out <= 16'h0243;    16'd41579: out <= 16'h0373;
    16'd41580: out <= 16'h0DF2;    16'd41581: out <= 16'h01F8;    16'd41582: out <= 16'h0811;    16'd41583: out <= 16'h068B;
    16'd41584: out <= 16'h017A;    16'd41585: out <= 16'h0636;    16'd41586: out <= 16'h04B6;    16'd41587: out <= 16'h0498;
    16'd41588: out <= 16'h0AB2;    16'd41589: out <= 16'h06F1;    16'd41590: out <= 16'h0323;    16'd41591: out <= 16'h053E;
    16'd41592: out <= 16'h06BC;    16'd41593: out <= 16'h0229;    16'd41594: out <= 16'h096D;    16'd41595: out <= 16'h0777;
    16'd41596: out <= 16'hFFA4;    16'd41597: out <= 16'hFD7D;    16'd41598: out <= 16'h00C5;    16'd41599: out <= 16'hFBF5;
    16'd41600: out <= 16'h0173;    16'd41601: out <= 16'h034C;    16'd41602: out <= 16'h02BB;    16'd41603: out <= 16'h0C03;
    16'd41604: out <= 16'h01F7;    16'd41605: out <= 16'h03A3;    16'd41606: out <= 16'h065C;    16'd41607: out <= 16'hFFB1;
    16'd41608: out <= 16'h063B;    16'd41609: out <= 16'h0788;    16'd41610: out <= 16'h065A;    16'd41611: out <= 16'h04B1;
    16'd41612: out <= 16'h02B7;    16'd41613: out <= 16'h0108;    16'd41614: out <= 16'h0285;    16'd41615: out <= 16'h0645;
    16'd41616: out <= 16'h0861;    16'd41617: out <= 16'h0516;    16'd41618: out <= 16'h00CD;    16'd41619: out <= 16'h0395;
    16'd41620: out <= 16'h040C;    16'd41621: out <= 16'h005B;    16'd41622: out <= 16'h0087;    16'd41623: out <= 16'h035C;
    16'd41624: out <= 16'hFE9C;    16'd41625: out <= 16'h0751;    16'd41626: out <= 16'h0363;    16'd41627: out <= 16'h048A;
    16'd41628: out <= 16'h00C9;    16'd41629: out <= 16'h03C2;    16'd41630: out <= 16'h0427;    16'd41631: out <= 16'h0276;
    16'd41632: out <= 16'h006C;    16'd41633: out <= 16'h0240;    16'd41634: out <= 16'hFD83;    16'd41635: out <= 16'h0A82;
    16'd41636: out <= 16'h0223;    16'd41637: out <= 16'h0591;    16'd41638: out <= 16'hFB80;    16'd41639: out <= 16'h025F;
    16'd41640: out <= 16'h07F5;    16'd41641: out <= 16'h0A04;    16'd41642: out <= 16'h03C7;    16'd41643: out <= 16'h03E2;
    16'd41644: out <= 16'h08ED;    16'd41645: out <= 16'h01B9;    16'd41646: out <= 16'h00B6;    16'd41647: out <= 16'h05F9;
    16'd41648: out <= 16'h04EE;    16'd41649: out <= 16'h06A2;    16'd41650: out <= 16'h0446;    16'd41651: out <= 16'h05DE;
    16'd41652: out <= 16'h0682;    16'd41653: out <= 16'h06A7;    16'd41654: out <= 16'h021B;    16'd41655: out <= 16'h01C9;
    16'd41656: out <= 16'h09D0;    16'd41657: out <= 16'h0144;    16'd41658: out <= 16'h04CC;    16'd41659: out <= 16'hFF16;
    16'd41660: out <= 16'h05FA;    16'd41661: out <= 16'hFE4D;    16'd41662: out <= 16'h010A;    16'd41663: out <= 16'h0AB1;
    16'd41664: out <= 16'h041A;    16'd41665: out <= 16'hFBC0;    16'd41666: out <= 16'h05AF;    16'd41667: out <= 16'h07A7;
    16'd41668: out <= 16'h08D4;    16'd41669: out <= 16'h0A92;    16'd41670: out <= 16'h0365;    16'd41671: out <= 16'h0795;
    16'd41672: out <= 16'h07CA;    16'd41673: out <= 16'hFF3B;    16'd41674: out <= 16'h0860;    16'd41675: out <= 16'h07B6;
    16'd41676: out <= 16'h0242;    16'd41677: out <= 16'h04DD;    16'd41678: out <= 16'h04D2;    16'd41679: out <= 16'h03C5;
    16'd41680: out <= 16'h022B;    16'd41681: out <= 16'h04F0;    16'd41682: out <= 16'h0601;    16'd41683: out <= 16'h07B1;
    16'd41684: out <= 16'h0A4B;    16'd41685: out <= 16'h03FB;    16'd41686: out <= 16'h02E2;    16'd41687: out <= 16'h05C5;
    16'd41688: out <= 16'h065C;    16'd41689: out <= 16'hFF41;    16'd41690: out <= 16'h0D03;    16'd41691: out <= 16'h0797;
    16'd41692: out <= 16'h0AD2;    16'd41693: out <= 16'h09B4;    16'd41694: out <= 16'h03A9;    16'd41695: out <= 16'h086E;
    16'd41696: out <= 16'hF727;    16'd41697: out <= 16'h01D2;    16'd41698: out <= 16'hFE4D;    16'd41699: out <= 16'h03A1;
    16'd41700: out <= 16'h00CF;    16'd41701: out <= 16'h01BC;    16'd41702: out <= 16'hFEEE;    16'd41703: out <= 16'h04B4;
    16'd41704: out <= 16'h0006;    16'd41705: out <= 16'h01D3;    16'd41706: out <= 16'hFA9C;    16'd41707: out <= 16'hFEE6;
    16'd41708: out <= 16'hF792;    16'd41709: out <= 16'h0542;    16'd41710: out <= 16'h03A8;    16'd41711: out <= 16'h0040;
    16'd41712: out <= 16'hFA52;    16'd41713: out <= 16'h01D2;    16'd41714: out <= 16'h0784;    16'd41715: out <= 16'h043D;
    16'd41716: out <= 16'h0380;    16'd41717: out <= 16'hFE02;    16'd41718: out <= 16'h0271;    16'd41719: out <= 16'h02CD;
    16'd41720: out <= 16'hFF58;    16'd41721: out <= 16'hFB90;    16'd41722: out <= 16'h012F;    16'd41723: out <= 16'hF9F3;
    16'd41724: out <= 16'h00A5;    16'd41725: out <= 16'hFEA8;    16'd41726: out <= 16'h01B2;    16'd41727: out <= 16'hFF31;
    16'd41728: out <= 16'h018F;    16'd41729: out <= 16'h01CB;    16'd41730: out <= 16'hFEB6;    16'd41731: out <= 16'h0128;
    16'd41732: out <= 16'h04EB;    16'd41733: out <= 16'hFD45;    16'd41734: out <= 16'h045E;    16'd41735: out <= 16'h04B5;
    16'd41736: out <= 16'h034C;    16'd41737: out <= 16'hFE43;    16'd41738: out <= 16'hFFD4;    16'd41739: out <= 16'h00A5;
    16'd41740: out <= 16'hFD79;    16'd41741: out <= 16'h0038;    16'd41742: out <= 16'hFF73;    16'd41743: out <= 16'hFC33;
    16'd41744: out <= 16'h0115;    16'd41745: out <= 16'hFBCB;    16'd41746: out <= 16'hFAF4;    16'd41747: out <= 16'h06A7;
    16'd41748: out <= 16'hFF42;    16'd41749: out <= 16'hFCFB;    16'd41750: out <= 16'hFDF3;    16'd41751: out <= 16'hFFA8;
    16'd41752: out <= 16'h0635;    16'd41753: out <= 16'h067F;    16'd41754: out <= 16'h02BD;    16'd41755: out <= 16'hF98E;
    16'd41756: out <= 16'hF9C2;    16'd41757: out <= 16'h0209;    16'd41758: out <= 16'h050D;    16'd41759: out <= 16'h0415;
    16'd41760: out <= 16'h044B;    16'd41761: out <= 16'h03AB;    16'd41762: out <= 16'h04DB;    16'd41763: out <= 16'hFF8C;
    16'd41764: out <= 16'h0412;    16'd41765: out <= 16'h00CB;    16'd41766: out <= 16'h065D;    16'd41767: out <= 16'h0AAD;
    16'd41768: out <= 16'h0761;    16'd41769: out <= 16'h08E7;    16'd41770: out <= 16'h03D5;    16'd41771: out <= 16'h0152;
    16'd41772: out <= 16'h0263;    16'd41773: out <= 16'hFFFF;    16'd41774: out <= 16'h030E;    16'd41775: out <= 16'h079A;
    16'd41776: out <= 16'h0712;    16'd41777: out <= 16'h079A;    16'd41778: out <= 16'h072D;    16'd41779: out <= 16'h06AA;
    16'd41780: out <= 16'h095E;    16'd41781: out <= 16'h036D;    16'd41782: out <= 16'h0503;    16'd41783: out <= 16'h07C4;
    16'd41784: out <= 16'h03A2;    16'd41785: out <= 16'h05DD;    16'd41786: out <= 16'h039D;    16'd41787: out <= 16'h076F;
    16'd41788: out <= 16'h0024;    16'd41789: out <= 16'h0406;    16'd41790: out <= 16'h04DC;    16'd41791: out <= 16'h0009;
    16'd41792: out <= 16'hFFEF;    16'd41793: out <= 16'h022E;    16'd41794: out <= 16'hFEAA;    16'd41795: out <= 16'h031E;
    16'd41796: out <= 16'hFAE1;    16'd41797: out <= 16'h0079;    16'd41798: out <= 16'h0C01;    16'd41799: out <= 16'h00E3;
    16'd41800: out <= 16'hFD03;    16'd41801: out <= 16'h0079;    16'd41802: out <= 16'h085B;    16'd41803: out <= 16'h03C3;
    16'd41804: out <= 16'h0A41;    16'd41805: out <= 16'h018C;    16'd41806: out <= 16'h04A2;    16'd41807: out <= 16'h0009;
    16'd41808: out <= 16'h032D;    16'd41809: out <= 16'h0C3C;    16'd41810: out <= 16'h0383;    16'd41811: out <= 16'h03D6;
    16'd41812: out <= 16'h0703;    16'd41813: out <= 16'h059B;    16'd41814: out <= 16'hFF07;    16'd41815: out <= 16'hFDB0;
    16'd41816: out <= 16'hFFE0;    16'd41817: out <= 16'h01C5;    16'd41818: out <= 16'h0023;    16'd41819: out <= 16'h0105;
    16'd41820: out <= 16'hFEE8;    16'd41821: out <= 16'h0656;    16'd41822: out <= 16'h05E8;    16'd41823: out <= 16'hFF52;
    16'd41824: out <= 16'h0496;    16'd41825: out <= 16'h0B07;    16'd41826: out <= 16'h01DA;    16'd41827: out <= 16'h0643;
    16'd41828: out <= 16'h02C4;    16'd41829: out <= 16'h007D;    16'd41830: out <= 16'h0840;    16'd41831: out <= 16'h070E;
    16'd41832: out <= 16'h07E1;    16'd41833: out <= 16'h0202;    16'd41834: out <= 16'h026D;    16'd41835: out <= 16'h0821;
    16'd41836: out <= 16'h07AA;    16'd41837: out <= 16'h0075;    16'd41838: out <= 16'h003E;    16'd41839: out <= 16'h0967;
    16'd41840: out <= 16'h00E2;    16'd41841: out <= 16'h0BEE;    16'd41842: out <= 16'h07FA;    16'd41843: out <= 16'h0578;
    16'd41844: out <= 16'h0194;    16'd41845: out <= 16'h025F;    16'd41846: out <= 16'h0203;    16'd41847: out <= 16'h0694;
    16'd41848: out <= 16'h071B;    16'd41849: out <= 16'h015C;    16'd41850: out <= 16'h042A;    16'd41851: out <= 16'hFF43;
    16'd41852: out <= 16'h07CA;    16'd41853: out <= 16'h058C;    16'd41854: out <= 16'hFCFF;    16'd41855: out <= 16'h03A3;
    16'd41856: out <= 16'h01E2;    16'd41857: out <= 16'h0845;    16'd41858: out <= 16'h0B2A;    16'd41859: out <= 16'h05A3;
    16'd41860: out <= 16'h0D96;    16'd41861: out <= 16'hFF7B;    16'd41862: out <= 16'h030F;    16'd41863: out <= 16'h08D5;
    16'd41864: out <= 16'h0649;    16'd41865: out <= 16'h05AD;    16'd41866: out <= 16'h0700;    16'd41867: out <= 16'h0465;
    16'd41868: out <= 16'h025B;    16'd41869: out <= 16'h0469;    16'd41870: out <= 16'hFE36;    16'd41871: out <= 16'h002F;
    16'd41872: out <= 16'h029E;    16'd41873: out <= 16'h036A;    16'd41874: out <= 16'h0464;    16'd41875: out <= 16'hFCA3;
    16'd41876: out <= 16'h0369;    16'd41877: out <= 16'h0452;    16'd41878: out <= 16'h0799;    16'd41879: out <= 16'h048D;
    16'd41880: out <= 16'h04DA;    16'd41881: out <= 16'h0097;    16'd41882: out <= 16'h029B;    16'd41883: out <= 16'h067A;
    16'd41884: out <= 16'h0252;    16'd41885: out <= 16'h0085;    16'd41886: out <= 16'h01BB;    16'd41887: out <= 16'h05E0;
    16'd41888: out <= 16'h0183;    16'd41889: out <= 16'h024B;    16'd41890: out <= 16'h0601;    16'd41891: out <= 16'h047E;
    16'd41892: out <= 16'h030F;    16'd41893: out <= 16'hFE33;    16'd41894: out <= 16'h02D9;    16'd41895: out <= 16'h089E;
    16'd41896: out <= 16'h02A3;    16'd41897: out <= 16'h08A2;    16'd41898: out <= 16'h0371;    16'd41899: out <= 16'h004A;
    16'd41900: out <= 16'h01F4;    16'd41901: out <= 16'h045B;    16'd41902: out <= 16'h01F1;    16'd41903: out <= 16'h0217;
    16'd41904: out <= 16'h05BB;    16'd41905: out <= 16'h00D2;    16'd41906: out <= 16'h0394;    16'd41907: out <= 16'h0842;
    16'd41908: out <= 16'h01C0;    16'd41909: out <= 16'h037B;    16'd41910: out <= 16'h0D60;    16'd41911: out <= 16'h08EA;
    16'd41912: out <= 16'h017D;    16'd41913: out <= 16'hFF1C;    16'd41914: out <= 16'h099D;    16'd41915: out <= 16'h02DC;
    16'd41916: out <= 16'h0639;    16'd41917: out <= 16'h0161;    16'd41918: out <= 16'h07F2;    16'd41919: out <= 16'h02A4;
    16'd41920: out <= 16'h06D1;    16'd41921: out <= 16'hFE71;    16'd41922: out <= 16'h08E3;    16'd41923: out <= 16'h075E;
    16'd41924: out <= 16'h08F3;    16'd41925: out <= 16'h019F;    16'd41926: out <= 16'h04AC;    16'd41927: out <= 16'h094A;
    16'd41928: out <= 16'hFEF3;    16'd41929: out <= 16'h0678;    16'd41930: out <= 16'h07A2;    16'd41931: out <= 16'h00D2;
    16'd41932: out <= 16'hFEBF;    16'd41933: out <= 16'h0329;    16'd41934: out <= 16'h0253;    16'd41935: out <= 16'h01DC;
    16'd41936: out <= 16'h03D4;    16'd41937: out <= 16'hFF32;    16'd41938: out <= 16'hFCB6;    16'd41939: out <= 16'h063A;
    16'd41940: out <= 16'h04C4;    16'd41941: out <= 16'h05D7;    16'd41942: out <= 16'h045D;    16'd41943: out <= 16'h0098;
    16'd41944: out <= 16'h0049;    16'd41945: out <= 16'h0342;    16'd41946: out <= 16'h02F4;    16'd41947: out <= 16'h0177;
    16'd41948: out <= 16'h0A7A;    16'd41949: out <= 16'h0A07;    16'd41950: out <= 16'h06A6;    16'd41951: out <= 16'h0102;
    16'd41952: out <= 16'hF9CA;    16'd41953: out <= 16'h0409;    16'd41954: out <= 16'h0C52;    16'd41955: out <= 16'hF7B8;
    16'd41956: out <= 16'hFDE8;    16'd41957: out <= 16'hFBB1;    16'd41958: out <= 16'h0069;    16'd41959: out <= 16'h0572;
    16'd41960: out <= 16'hFE64;    16'd41961: out <= 16'hFFC0;    16'd41962: out <= 16'h00A7;    16'd41963: out <= 16'h0315;
    16'd41964: out <= 16'h041A;    16'd41965: out <= 16'h01C1;    16'd41966: out <= 16'hFDAC;    16'd41967: out <= 16'h059B;
    16'd41968: out <= 16'h0134;    16'd41969: out <= 16'h00E9;    16'd41970: out <= 16'h00D6;    16'd41971: out <= 16'hFD7B;
    16'd41972: out <= 16'hFD1A;    16'd41973: out <= 16'h01E4;    16'd41974: out <= 16'h032C;    16'd41975: out <= 16'hFF5D;
    16'd41976: out <= 16'hFB7F;    16'd41977: out <= 16'h03A9;    16'd41978: out <= 16'hFDEA;    16'd41979: out <= 16'h0636;
    16'd41980: out <= 16'hF76D;    16'd41981: out <= 16'h0606;    16'd41982: out <= 16'h013F;    16'd41983: out <= 16'hFFAB;
    16'd41984: out <= 16'h0252;    16'd41985: out <= 16'hFEA0;    16'd41986: out <= 16'hFFC1;    16'd41987: out <= 16'hFCAB;
    16'd41988: out <= 16'hFD87;    16'd41989: out <= 16'h02AD;    16'd41990: out <= 16'h00C3;    16'd41991: out <= 16'hFCA8;
    16'd41992: out <= 16'h02EB;    16'd41993: out <= 16'h034B;    16'd41994: out <= 16'hFD91;    16'd41995: out <= 16'h063D;
    16'd41996: out <= 16'hF874;    16'd41997: out <= 16'hFF27;    16'd41998: out <= 16'h037F;    16'd41999: out <= 16'hFC00;
    16'd42000: out <= 16'hFD7F;    16'd42001: out <= 16'h09E0;    16'd42002: out <= 16'h01F1;    16'd42003: out <= 16'hFE0E;
    16'd42004: out <= 16'h009F;    16'd42005: out <= 16'hFFBB;    16'd42006: out <= 16'h0224;    16'd42007: out <= 16'h02A5;
    16'd42008: out <= 16'h030F;    16'd42009: out <= 16'h0492;    16'd42010: out <= 16'h01A4;    16'd42011: out <= 16'hFB7B;
    16'd42012: out <= 16'hFFE0;    16'd42013: out <= 16'hFA90;    16'd42014: out <= 16'h01D4;    16'd42015: out <= 16'h0528;
    16'd42016: out <= 16'h04B6;    16'd42017: out <= 16'h05C2;    16'd42018: out <= 16'hFE13;    16'd42019: out <= 16'h02B0;
    16'd42020: out <= 16'h0394;    16'd42021: out <= 16'h0336;    16'd42022: out <= 16'h0953;    16'd42023: out <= 16'h0298;
    16'd42024: out <= 16'hFC5F;    16'd42025: out <= 16'h01F0;    16'd42026: out <= 16'h015E;    16'd42027: out <= 16'h032F;
    16'd42028: out <= 16'h0949;    16'd42029: out <= 16'h04EB;    16'd42030: out <= 16'h03A1;    16'd42031: out <= 16'h08AD;
    16'd42032: out <= 16'h0382;    16'd42033: out <= 16'h0449;    16'd42034: out <= 16'h05A7;    16'd42035: out <= 16'h0031;
    16'd42036: out <= 16'h062E;    16'd42037: out <= 16'h032B;    16'd42038: out <= 16'hFFC4;    16'd42039: out <= 16'h0A5F;
    16'd42040: out <= 16'h0806;    16'd42041: out <= 16'hFB87;    16'd42042: out <= 16'hFF9F;    16'd42043: out <= 16'h0C9D;
    16'd42044: out <= 16'h027E;    16'd42045: out <= 16'h0C77;    16'd42046: out <= 16'h0705;    16'd42047: out <= 16'h0016;
    16'd42048: out <= 16'h0A84;    16'd42049: out <= 16'hFF70;    16'd42050: out <= 16'h01FD;    16'd42051: out <= 16'h0272;
    16'd42052: out <= 16'hFE4F;    16'd42053: out <= 16'hFD53;    16'd42054: out <= 16'h02A6;    16'd42055: out <= 16'h0165;
    16'd42056: out <= 16'h06C2;    16'd42057: out <= 16'h05D4;    16'd42058: out <= 16'h0664;    16'd42059: out <= 16'h058F;
    16'd42060: out <= 16'h043B;    16'd42061: out <= 16'h02B5;    16'd42062: out <= 16'h0422;    16'd42063: out <= 16'h01B6;
    16'd42064: out <= 16'h065D;    16'd42065: out <= 16'h0834;    16'd42066: out <= 16'hFB97;    16'd42067: out <= 16'h039C;
    16'd42068: out <= 16'h0449;    16'd42069: out <= 16'h0461;    16'd42070: out <= 16'h052B;    16'd42071: out <= 16'h0418;
    16'd42072: out <= 16'h03E1;    16'd42073: out <= 16'hFCAE;    16'd42074: out <= 16'h006E;    16'd42075: out <= 16'h008C;
    16'd42076: out <= 16'h075D;    16'd42077: out <= 16'hFF1D;    16'd42078: out <= 16'h0765;    16'd42079: out <= 16'h026F;
    16'd42080: out <= 16'h07B6;    16'd42081: out <= 16'h0495;    16'd42082: out <= 16'h0743;    16'd42083: out <= 16'h0670;
    16'd42084: out <= 16'h0068;    16'd42085: out <= 16'h00F8;    16'd42086: out <= 16'h0023;    16'd42087: out <= 16'h0287;
    16'd42088: out <= 16'hFC6B;    16'd42089: out <= 16'h0609;    16'd42090: out <= 16'hFE62;    16'd42091: out <= 16'h01DD;
    16'd42092: out <= 16'h03F4;    16'd42093: out <= 16'h076E;    16'd42094: out <= 16'h061E;    16'd42095: out <= 16'h07B0;
    16'd42096: out <= 16'h020D;    16'd42097: out <= 16'h07D3;    16'd42098: out <= 16'h0622;    16'd42099: out <= 16'h02CF;
    16'd42100: out <= 16'h0392;    16'd42101: out <= 16'h0647;    16'd42102: out <= 16'h0395;    16'd42103: out <= 16'h06E0;
    16'd42104: out <= 16'h00E9;    16'd42105: out <= 16'h04DA;    16'd42106: out <= 16'h079F;    16'd42107: out <= 16'h020B;
    16'd42108: out <= 16'hFC31;    16'd42109: out <= 16'h05AB;    16'd42110: out <= 16'h0521;    16'd42111: out <= 16'h0712;
    16'd42112: out <= 16'h09D2;    16'd42113: out <= 16'h0094;    16'd42114: out <= 16'hF94D;    16'd42115: out <= 16'h0598;
    16'd42116: out <= 16'h0016;    16'd42117: out <= 16'h044C;    16'd42118: out <= 16'h001B;    16'd42119: out <= 16'h000C;
    16'd42120: out <= 16'h05AA;    16'd42121: out <= 16'h04DA;    16'd42122: out <= 16'h09B9;    16'd42123: out <= 16'h020A;
    16'd42124: out <= 16'h080B;    16'd42125: out <= 16'hFBFE;    16'd42126: out <= 16'h05E2;    16'd42127: out <= 16'h0686;
    16'd42128: out <= 16'h059B;    16'd42129: out <= 16'h04F9;    16'd42130: out <= 16'h0610;    16'd42131: out <= 16'h0867;
    16'd42132: out <= 16'h01BE;    16'd42133: out <= 16'h05DF;    16'd42134: out <= 16'h01D7;    16'd42135: out <= 16'hFE34;
    16'd42136: out <= 16'hFF65;    16'd42137: out <= 16'h07F8;    16'd42138: out <= 16'hFF65;    16'd42139: out <= 16'h0723;
    16'd42140: out <= 16'h02B3;    16'd42141: out <= 16'h059B;    16'd42142: out <= 16'h058A;    16'd42143: out <= 16'h0940;
    16'd42144: out <= 16'h0C2B;    16'd42145: out <= 16'h0474;    16'd42146: out <= 16'hFD15;    16'd42147: out <= 16'h067C;
    16'd42148: out <= 16'h0481;    16'd42149: out <= 16'h07E9;    16'd42150: out <= 16'h0385;    16'd42151: out <= 16'h0276;
    16'd42152: out <= 16'h0691;    16'd42153: out <= 16'h0407;    16'd42154: out <= 16'h051B;    16'd42155: out <= 16'h022F;
    16'd42156: out <= 16'h01A4;    16'd42157: out <= 16'h04E3;    16'd42158: out <= 16'h0283;    16'd42159: out <= 16'h0258;
    16'd42160: out <= 16'h0882;    16'd42161: out <= 16'h08C5;    16'd42162: out <= 16'h0301;    16'd42163: out <= 16'h08BF;
    16'd42164: out <= 16'hFB03;    16'd42165: out <= 16'h03D6;    16'd42166: out <= 16'hFFD1;    16'd42167: out <= 16'hFABC;
    16'd42168: out <= 16'h02C9;    16'd42169: out <= 16'h038D;    16'd42170: out <= 16'h0532;    16'd42171: out <= 16'h028F;
    16'd42172: out <= 16'hFDE8;    16'd42173: out <= 16'h02C7;    16'd42174: out <= 16'h086F;    16'd42175: out <= 16'h069A;
    16'd42176: out <= 16'h08ED;    16'd42177: out <= 16'h0402;    16'd42178: out <= 16'h0B29;    16'd42179: out <= 16'h0800;
    16'd42180: out <= 16'h0252;    16'd42181: out <= 16'h03A8;    16'd42182: out <= 16'h01F6;    16'd42183: out <= 16'h039D;
    16'd42184: out <= 16'h0258;    16'd42185: out <= 16'h059D;    16'd42186: out <= 16'h03AD;    16'd42187: out <= 16'hFF4A;
    16'd42188: out <= 16'h030B;    16'd42189: out <= 16'h024F;    16'd42190: out <= 16'hFCA6;    16'd42191: out <= 16'h088A;
    16'd42192: out <= 16'h0516;    16'd42193: out <= 16'h0124;    16'd42194: out <= 16'h0733;    16'd42195: out <= 16'h02AA;
    16'd42196: out <= 16'h062F;    16'd42197: out <= 16'h08F1;    16'd42198: out <= 16'h023F;    16'd42199: out <= 16'h0101;
    16'd42200: out <= 16'h03EF;    16'd42201: out <= 16'h013B;    16'd42202: out <= 16'h039C;    16'd42203: out <= 16'h04ED;
    16'd42204: out <= 16'h01FA;    16'd42205: out <= 16'hFC6D;    16'd42206: out <= 16'h0567;    16'd42207: out <= 16'h05E7;
    16'd42208: out <= 16'hFD38;    16'd42209: out <= 16'h00F4;    16'd42210: out <= 16'hFCB8;    16'd42211: out <= 16'hFF94;
    16'd42212: out <= 16'h0666;    16'd42213: out <= 16'h00E3;    16'd42214: out <= 16'hFC42;    16'd42215: out <= 16'hFF6C;
    16'd42216: out <= 16'h03C3;    16'd42217: out <= 16'hFF72;    16'd42218: out <= 16'hFC92;    16'd42219: out <= 16'hFD4A;
    16'd42220: out <= 16'hFBE0;    16'd42221: out <= 16'hF9B2;    16'd42222: out <= 16'hFF9F;    16'd42223: out <= 16'hFEC1;
    16'd42224: out <= 16'h037B;    16'd42225: out <= 16'hFE3E;    16'd42226: out <= 16'h021D;    16'd42227: out <= 16'hFD1A;
    16'd42228: out <= 16'h0188;    16'd42229: out <= 16'hF908;    16'd42230: out <= 16'hFD6E;    16'd42231: out <= 16'hFF46;
    16'd42232: out <= 16'h02DA;    16'd42233: out <= 16'hFE33;    16'd42234: out <= 16'hFB4F;    16'd42235: out <= 16'hFACF;
    16'd42236: out <= 16'hFBCE;    16'd42237: out <= 16'hFE54;    16'd42238: out <= 16'hFED1;    16'd42239: out <= 16'hFE71;
    16'd42240: out <= 16'h08D7;    16'd42241: out <= 16'hFCF2;    16'd42242: out <= 16'hFE1B;    16'd42243: out <= 16'h03FA;
    16'd42244: out <= 16'h00E8;    16'd42245: out <= 16'h0753;    16'd42246: out <= 16'h0357;    16'd42247: out <= 16'hFAA0;
    16'd42248: out <= 16'h0411;    16'd42249: out <= 16'h00D1;    16'd42250: out <= 16'hFE2D;    16'd42251: out <= 16'h007C;
    16'd42252: out <= 16'h0200;    16'd42253: out <= 16'h0370;    16'd42254: out <= 16'hFCB2;    16'd42255: out <= 16'h0155;
    16'd42256: out <= 16'h04FF;    16'd42257: out <= 16'hFDDB;    16'd42258: out <= 16'hFDF6;    16'd42259: out <= 16'hF71E;
    16'd42260: out <= 16'hFFD5;    16'd42261: out <= 16'h005F;    16'd42262: out <= 16'hFAAD;    16'd42263: out <= 16'h036D;
    16'd42264: out <= 16'hF965;    16'd42265: out <= 16'hFB60;    16'd42266: out <= 16'hFF32;    16'd42267: out <= 16'h0134;
    16'd42268: out <= 16'hFC14;    16'd42269: out <= 16'hFE8A;    16'd42270: out <= 16'h0113;    16'd42271: out <= 16'hFFAF;
    16'd42272: out <= 16'h04B0;    16'd42273: out <= 16'h008E;    16'd42274: out <= 16'hFF25;    16'd42275: out <= 16'h04E5;
    16'd42276: out <= 16'h0857;    16'd42277: out <= 16'h032B;    16'd42278: out <= 16'h01E4;    16'd42279: out <= 16'h039D;
    16'd42280: out <= 16'h0110;    16'd42281: out <= 16'h079C;    16'd42282: out <= 16'h05FB;    16'd42283: out <= 16'h03D2;
    16'd42284: out <= 16'h08EA;    16'd42285: out <= 16'h0785;    16'd42286: out <= 16'h05CE;    16'd42287: out <= 16'h07C1;
    16'd42288: out <= 16'h044C;    16'd42289: out <= 16'hFEED;    16'd42290: out <= 16'h02A3;    16'd42291: out <= 16'h05EB;
    16'd42292: out <= 16'h091D;    16'd42293: out <= 16'h04D1;    16'd42294: out <= 16'h035C;    16'd42295: out <= 16'h040E;
    16'd42296: out <= 16'h03D7;    16'd42297: out <= 16'hFF95;    16'd42298: out <= 16'h036F;    16'd42299: out <= 16'hFF2D;
    16'd42300: out <= 16'hFF95;    16'd42301: out <= 16'h09FE;    16'd42302: out <= 16'h04D9;    16'd42303: out <= 16'h07DE;
    16'd42304: out <= 16'h0905;    16'd42305: out <= 16'h0428;    16'd42306: out <= 16'h0721;    16'd42307: out <= 16'h05C8;
    16'd42308: out <= 16'h0645;    16'd42309: out <= 16'hFD8D;    16'd42310: out <= 16'h0AD8;    16'd42311: out <= 16'h0BEF;
    16'd42312: out <= 16'h0309;    16'd42313: out <= 16'h00EF;    16'd42314: out <= 16'h0860;    16'd42315: out <= 16'h0432;
    16'd42316: out <= 16'h0549;    16'd42317: out <= 16'h02B5;    16'd42318: out <= 16'h0317;    16'd42319: out <= 16'h0A6C;
    16'd42320: out <= 16'h0699;    16'd42321: out <= 16'hFFDF;    16'd42322: out <= 16'hFF90;    16'd42323: out <= 16'h0228;
    16'd42324: out <= 16'h0740;    16'd42325: out <= 16'h0596;    16'd42326: out <= 16'hFF04;    16'd42327: out <= 16'h074A;
    16'd42328: out <= 16'h02B7;    16'd42329: out <= 16'h0649;    16'd42330: out <= 16'h0489;    16'd42331: out <= 16'hFC87;
    16'd42332: out <= 16'h0079;    16'd42333: out <= 16'h0480;    16'd42334: out <= 16'h0270;    16'd42335: out <= 16'hFE8A;
    16'd42336: out <= 16'h092C;    16'd42337: out <= 16'h0290;    16'd42338: out <= 16'h0083;    16'd42339: out <= 16'hFF89;
    16'd42340: out <= 16'h0BED;    16'd42341: out <= 16'h0480;    16'd42342: out <= 16'hFF1E;    16'd42343: out <= 16'h05E5;
    16'd42344: out <= 16'hFC97;    16'd42345: out <= 16'hFCA8;    16'd42346: out <= 16'hFF78;    16'd42347: out <= 16'h076E;
    16'd42348: out <= 16'h005D;    16'd42349: out <= 16'h03CA;    16'd42350: out <= 16'h0740;    16'd42351: out <= 16'h024C;
    16'd42352: out <= 16'h0366;    16'd42353: out <= 16'hFFC9;    16'd42354: out <= 16'h045C;    16'd42355: out <= 16'h0035;
    16'd42356: out <= 16'h05F5;    16'd42357: out <= 16'h03B7;    16'd42358: out <= 16'hFF7A;    16'd42359: out <= 16'h031E;
    16'd42360: out <= 16'h0AB9;    16'd42361: out <= 16'h0255;    16'd42362: out <= 16'h0538;    16'd42363: out <= 16'h0244;
    16'd42364: out <= 16'hFFC7;    16'd42365: out <= 16'h0834;    16'd42366: out <= 16'h02D6;    16'd42367: out <= 16'h0389;
    16'd42368: out <= 16'hFF38;    16'd42369: out <= 16'hFCDD;    16'd42370: out <= 16'h0587;    16'd42371: out <= 16'h0564;
    16'd42372: out <= 16'h05DF;    16'd42373: out <= 16'hFF1D;    16'd42374: out <= 16'h0201;    16'd42375: out <= 16'h0167;
    16'd42376: out <= 16'h02D8;    16'd42377: out <= 16'h06BC;    16'd42378: out <= 16'h08F3;    16'd42379: out <= 16'h0849;
    16'd42380: out <= 16'h0CFC;    16'd42381: out <= 16'h0562;    16'd42382: out <= 16'h0812;    16'd42383: out <= 16'h01D4;
    16'd42384: out <= 16'h0976;    16'd42385: out <= 16'h043E;    16'd42386: out <= 16'h0280;    16'd42387: out <= 16'h00C5;
    16'd42388: out <= 16'h0358;    16'd42389: out <= 16'h06D9;    16'd42390: out <= 16'h025F;    16'd42391: out <= 16'h0662;
    16'd42392: out <= 16'h04AA;    16'd42393: out <= 16'h068C;    16'd42394: out <= 16'h0687;    16'd42395: out <= 16'hFEDC;
    16'd42396: out <= 16'hFF1C;    16'd42397: out <= 16'h0A7B;    16'd42398: out <= 16'h0673;    16'd42399: out <= 16'h0A13;
    16'd42400: out <= 16'h0728;    16'd42401: out <= 16'h05CF;    16'd42402: out <= 16'hFFE8;    16'd42403: out <= 16'hFFDE;
    16'd42404: out <= 16'h0328;    16'd42405: out <= 16'h0B1D;    16'd42406: out <= 16'h0311;    16'd42407: out <= 16'h0A87;
    16'd42408: out <= 16'hFFE0;    16'd42409: out <= 16'h0573;    16'd42410: out <= 16'h0448;    16'd42411: out <= 16'h04A2;
    16'd42412: out <= 16'h00EB;    16'd42413: out <= 16'hFE6B;    16'd42414: out <= 16'hFE97;    16'd42415: out <= 16'h0EF5;
    16'd42416: out <= 16'h02EE;    16'd42417: out <= 16'h01D2;    16'd42418: out <= 16'h01FD;    16'd42419: out <= 16'h09A9;
    16'd42420: out <= 16'h0860;    16'd42421: out <= 16'h0032;    16'd42422: out <= 16'h069D;    16'd42423: out <= 16'h04C0;
    16'd42424: out <= 16'h01BC;    16'd42425: out <= 16'h0884;    16'd42426: out <= 16'h059A;    16'd42427: out <= 16'hFE63;
    16'd42428: out <= 16'h0384;    16'd42429: out <= 16'hFE41;    16'd42430: out <= 16'hFAF2;    16'd42431: out <= 16'hFF13;
    16'd42432: out <= 16'hFD76;    16'd42433: out <= 16'h01A2;    16'd42434: out <= 16'h064A;    16'd42435: out <= 16'hFFD8;
    16'd42436: out <= 16'hFEDD;    16'd42437: out <= 16'h066F;    16'd42438: out <= 16'h0801;    16'd42439: out <= 16'h01F1;
    16'd42440: out <= 16'h03DE;    16'd42441: out <= 16'h0280;    16'd42442: out <= 16'h0388;    16'd42443: out <= 16'h0295;
    16'd42444: out <= 16'h01AC;    16'd42445: out <= 16'h037E;    16'd42446: out <= 16'h04B7;    16'd42447: out <= 16'h0B16;
    16'd42448: out <= 16'h054D;    16'd42449: out <= 16'hFAA6;    16'd42450: out <= 16'h0439;    16'd42451: out <= 16'h0449;
    16'd42452: out <= 16'h008D;    16'd42453: out <= 16'h0865;    16'd42454: out <= 16'h0624;    16'd42455: out <= 16'h08AC;
    16'd42456: out <= 16'h0B7A;    16'd42457: out <= 16'h08FC;    16'd42458: out <= 16'h03F4;    16'd42459: out <= 16'h0A7D;
    16'd42460: out <= 16'h027F;    16'd42461: out <= 16'h087F;    16'd42462: out <= 16'hFB1E;    16'd42463: out <= 16'hFFA3;
    16'd42464: out <= 16'h005D;    16'd42465: out <= 16'hFF9D;    16'd42466: out <= 16'hF30D;    16'd42467: out <= 16'h0596;
    16'd42468: out <= 16'h044A;    16'd42469: out <= 16'h01A6;    16'd42470: out <= 16'hFEDD;    16'd42471: out <= 16'h048F;
    16'd42472: out <= 16'hF889;    16'd42473: out <= 16'hFB0B;    16'd42474: out <= 16'hFD33;    16'd42475: out <= 16'h0433;
    16'd42476: out <= 16'hFD40;    16'd42477: out <= 16'hFB4F;    16'd42478: out <= 16'h0419;    16'd42479: out <= 16'hFF47;
    16'd42480: out <= 16'hFEE4;    16'd42481: out <= 16'h03B0;    16'd42482: out <= 16'h02F6;    16'd42483: out <= 16'hFF7C;
    16'd42484: out <= 16'h0368;    16'd42485: out <= 16'h023C;    16'd42486: out <= 16'h009C;    16'd42487: out <= 16'hFDEA;
    16'd42488: out <= 16'hF6E5;    16'd42489: out <= 16'hFBF8;    16'd42490: out <= 16'hFCB9;    16'd42491: out <= 16'h0781;
    16'd42492: out <= 16'hFA9E;    16'd42493: out <= 16'hFFA3;    16'd42494: out <= 16'h055E;    16'd42495: out <= 16'hF728;
    16'd42496: out <= 16'hFB77;    16'd42497: out <= 16'hFFE0;    16'd42498: out <= 16'h0595;    16'd42499: out <= 16'hFA74;
    16'd42500: out <= 16'hFEE4;    16'd42501: out <= 16'hFE3C;    16'd42502: out <= 16'h010C;    16'd42503: out <= 16'h00B6;
    16'd42504: out <= 16'h05AA;    16'd42505: out <= 16'hFAE5;    16'd42506: out <= 16'h079D;    16'd42507: out <= 16'hFFEA;
    16'd42508: out <= 16'h03AA;    16'd42509: out <= 16'h0311;    16'd42510: out <= 16'h05FE;    16'd42511: out <= 16'h01AF;
    16'd42512: out <= 16'hFC6C;    16'd42513: out <= 16'hF99F;    16'd42514: out <= 16'hFF03;    16'd42515: out <= 16'hFF7B;
    16'd42516: out <= 16'hFA59;    16'd42517: out <= 16'hFFC6;    16'd42518: out <= 16'hF8B3;    16'd42519: out <= 16'hFFEE;
    16'd42520: out <= 16'hFD98;    16'd42521: out <= 16'hFB24;    16'd42522: out <= 16'h0559;    16'd42523: out <= 16'h020F;
    16'd42524: out <= 16'hFDA9;    16'd42525: out <= 16'hFF94;    16'd42526: out <= 16'h013E;    16'd42527: out <= 16'h0A37;
    16'd42528: out <= 16'h05B9;    16'd42529: out <= 16'h0549;    16'd42530: out <= 16'h08F1;    16'd42531: out <= 16'h021C;
    16'd42532: out <= 16'h00C3;    16'd42533: out <= 16'h0620;    16'd42534: out <= 16'h085E;    16'd42535: out <= 16'h012E;
    16'd42536: out <= 16'h0836;    16'd42537: out <= 16'hF98E;    16'd42538: out <= 16'h0905;    16'd42539: out <= 16'h05CA;
    16'd42540: out <= 16'h0982;    16'd42541: out <= 16'h0636;    16'd42542: out <= 16'h0343;    16'd42543: out <= 16'h0D51;
    16'd42544: out <= 16'hFF77;    16'd42545: out <= 16'h078E;    16'd42546: out <= 16'h05F9;    16'd42547: out <= 16'h002D;
    16'd42548: out <= 16'h004A;    16'd42549: out <= 16'h019F;    16'd42550: out <= 16'h02FA;    16'd42551: out <= 16'h0318;
    16'd42552: out <= 16'h0515;    16'd42553: out <= 16'h0114;    16'd42554: out <= 16'h0A51;    16'd42555: out <= 16'h0818;
    16'd42556: out <= 16'h0231;    16'd42557: out <= 16'h06E7;    16'd42558: out <= 16'h076A;    16'd42559: out <= 16'hFE56;
    16'd42560: out <= 16'h03E9;    16'd42561: out <= 16'h06C0;    16'd42562: out <= 16'h03A9;    16'd42563: out <= 16'h03DB;
    16'd42564: out <= 16'h0582;    16'd42565: out <= 16'h05D9;    16'd42566: out <= 16'h07FD;    16'd42567: out <= 16'h044D;
    16'd42568: out <= 16'h0345;    16'd42569: out <= 16'h0999;    16'd42570: out <= 16'h0144;    16'd42571: out <= 16'h01DC;
    16'd42572: out <= 16'h02DB;    16'd42573: out <= 16'h0324;    16'd42574: out <= 16'hFC8D;    16'd42575: out <= 16'h0441;
    16'd42576: out <= 16'h05D8;    16'd42577: out <= 16'h05D4;    16'd42578: out <= 16'h0988;    16'd42579: out <= 16'h08B4;
    16'd42580: out <= 16'h0858;    16'd42581: out <= 16'hFF94;    16'd42582: out <= 16'h0071;    16'd42583: out <= 16'h07A4;
    16'd42584: out <= 16'h02D8;    16'd42585: out <= 16'h01E9;    16'd42586: out <= 16'hFFDB;    16'd42587: out <= 16'h0514;
    16'd42588: out <= 16'hFF26;    16'd42589: out <= 16'h070E;    16'd42590: out <= 16'hFE13;    16'd42591: out <= 16'h02AB;
    16'd42592: out <= 16'h07D9;    16'd42593: out <= 16'h0BAC;    16'd42594: out <= 16'h0423;    16'd42595: out <= 16'hFA98;
    16'd42596: out <= 16'h00FE;    16'd42597: out <= 16'hFF33;    16'd42598: out <= 16'h04CC;    16'd42599: out <= 16'h0480;
    16'd42600: out <= 16'hFC89;    16'd42601: out <= 16'h0F71;    16'd42602: out <= 16'hFE22;    16'd42603: out <= 16'hFD58;
    16'd42604: out <= 16'h04C9;    16'd42605: out <= 16'h03F7;    16'd42606: out <= 16'h05AC;    16'd42607: out <= 16'h02E9;
    16'd42608: out <= 16'h051A;    16'd42609: out <= 16'h07F6;    16'd42610: out <= 16'hFEA6;    16'd42611: out <= 16'h031B;
    16'd42612: out <= 16'h0A78;    16'd42613: out <= 16'h06C1;    16'd42614: out <= 16'h06E6;    16'd42615: out <= 16'h02F3;
    16'd42616: out <= 16'h0787;    16'd42617: out <= 16'h0765;    16'd42618: out <= 16'h0419;    16'd42619: out <= 16'h038D;
    16'd42620: out <= 16'h08DD;    16'd42621: out <= 16'h0675;    16'd42622: out <= 16'h0888;    16'd42623: out <= 16'h013F;
    16'd42624: out <= 16'h0479;    16'd42625: out <= 16'h07BF;    16'd42626: out <= 16'h016C;    16'd42627: out <= 16'h0659;
    16'd42628: out <= 16'h04BF;    16'd42629: out <= 16'h0511;    16'd42630: out <= 16'h0477;    16'd42631: out <= 16'h0217;
    16'd42632: out <= 16'hFE00;    16'd42633: out <= 16'h023E;    16'd42634: out <= 16'h0267;    16'd42635: out <= 16'h0310;
    16'd42636: out <= 16'h0435;    16'd42637: out <= 16'h0262;    16'd42638: out <= 16'hFF17;    16'd42639: out <= 16'h002A;
    16'd42640: out <= 16'h062A;    16'd42641: out <= 16'h02D9;    16'd42642: out <= 16'h079B;    16'd42643: out <= 16'h07F5;
    16'd42644: out <= 16'h075B;    16'd42645: out <= 16'h0501;    16'd42646: out <= 16'h04E3;    16'd42647: out <= 16'h0B20;
    16'd42648: out <= 16'h05D9;    16'd42649: out <= 16'h0383;    16'd42650: out <= 16'h081F;    16'd42651: out <= 16'h085E;
    16'd42652: out <= 16'h0207;    16'd42653: out <= 16'h062B;    16'd42654: out <= 16'h0447;    16'd42655: out <= 16'h0081;
    16'd42656: out <= 16'h03B5;    16'd42657: out <= 16'h026C;    16'd42658: out <= 16'h067F;    16'd42659: out <= 16'h0292;
    16'd42660: out <= 16'h024E;    16'd42661: out <= 16'h051B;    16'd42662: out <= 16'h0A5A;    16'd42663: out <= 16'hFD8A;
    16'd42664: out <= 16'h06F2;    16'd42665: out <= 16'hFE21;    16'd42666: out <= 16'h0044;    16'd42667: out <= 16'h00E3;
    16'd42668: out <= 16'h066D;    16'd42669: out <= 16'h0025;    16'd42670: out <= 16'h013F;    16'd42671: out <= 16'h067E;
    16'd42672: out <= 16'h0589;    16'd42673: out <= 16'h040E;    16'd42674: out <= 16'h0740;    16'd42675: out <= 16'h093C;
    16'd42676: out <= 16'h032B;    16'd42677: out <= 16'h062E;    16'd42678: out <= 16'h075A;    16'd42679: out <= 16'h02D3;
    16'd42680: out <= 16'h0237;    16'd42681: out <= 16'h08EF;    16'd42682: out <= 16'h02B9;    16'd42683: out <= 16'hFDB6;
    16'd42684: out <= 16'h05EA;    16'd42685: out <= 16'h0021;    16'd42686: out <= 16'hFF91;    16'd42687: out <= 16'h0209;
    16'd42688: out <= 16'h042A;    16'd42689: out <= 16'h0410;    16'd42690: out <= 16'h03FF;    16'd42691: out <= 16'h022D;
    16'd42692: out <= 16'hFCE1;    16'd42693: out <= 16'hFF78;    16'd42694: out <= 16'h0065;    16'd42695: out <= 16'h0386;
    16'd42696: out <= 16'h0952;    16'd42697: out <= 16'h0769;    16'd42698: out <= 16'h03D3;    16'd42699: out <= 16'h05CE;
    16'd42700: out <= 16'h01B2;    16'd42701: out <= 16'h04EC;    16'd42702: out <= 16'hFFBF;    16'd42703: out <= 16'h02BA;
    16'd42704: out <= 16'h0434;    16'd42705: out <= 16'hFF4B;    16'd42706: out <= 16'h0C1B;    16'd42707: out <= 16'h05A2;
    16'd42708: out <= 16'h0649;    16'd42709: out <= 16'h03AC;    16'd42710: out <= 16'hFAC1;    16'd42711: out <= 16'h00E1;
    16'd42712: out <= 16'h0368;    16'd42713: out <= 16'h03E4;    16'd42714: out <= 16'h03F5;    16'd42715: out <= 16'h018A;
    16'd42716: out <= 16'h0A77;    16'd42717: out <= 16'h012B;    16'd42718: out <= 16'h00CF;    16'd42719: out <= 16'hFB70;
    16'd42720: out <= 16'h01D3;    16'd42721: out <= 16'h0066;    16'd42722: out <= 16'h03E5;    16'd42723: out <= 16'h0527;
    16'd42724: out <= 16'hFCD5;    16'd42725: out <= 16'hFBC0;    16'd42726: out <= 16'h0101;    16'd42727: out <= 16'h0264;
    16'd42728: out <= 16'hFEF6;    16'd42729: out <= 16'h015C;    16'd42730: out <= 16'h00F8;    16'd42731: out <= 16'h02BA;
    16'd42732: out <= 16'h0010;    16'd42733: out <= 16'h036E;    16'd42734: out <= 16'h04DF;    16'd42735: out <= 16'hFA94;
    16'd42736: out <= 16'h019C;    16'd42737: out <= 16'h03E5;    16'd42738: out <= 16'h03A9;    16'd42739: out <= 16'hFDC5;
    16'd42740: out <= 16'hFD5A;    16'd42741: out <= 16'h07CD;    16'd42742: out <= 16'h02A4;    16'd42743: out <= 16'h012B;
    16'd42744: out <= 16'h0267;    16'd42745: out <= 16'h08AD;    16'd42746: out <= 16'hFCE6;    16'd42747: out <= 16'hFF6D;
    16'd42748: out <= 16'h04B1;    16'd42749: out <= 16'h046F;    16'd42750: out <= 16'h02F3;    16'd42751: out <= 16'hFFB5;
    16'd42752: out <= 16'hFE07;    16'd42753: out <= 16'hFFD3;    16'd42754: out <= 16'hFFAE;    16'd42755: out <= 16'hFDF0;
    16'd42756: out <= 16'hFF67;    16'd42757: out <= 16'h047E;    16'd42758: out <= 16'hFDB6;    16'd42759: out <= 16'h00B9;
    16'd42760: out <= 16'h01E4;    16'd42761: out <= 16'h0846;    16'd42762: out <= 16'hFFE4;    16'd42763: out <= 16'h0026;
    16'd42764: out <= 16'h02F8;    16'd42765: out <= 16'h00FD;    16'd42766: out <= 16'h01CA;    16'd42767: out <= 16'h0402;
    16'd42768: out <= 16'h0355;    16'd42769: out <= 16'h034A;    16'd42770: out <= 16'hFE79;    16'd42771: out <= 16'h0235;
    16'd42772: out <= 16'h035F;    16'd42773: out <= 16'hFCB0;    16'd42774: out <= 16'h004E;    16'd42775: out <= 16'hFFD5;
    16'd42776: out <= 16'h0463;    16'd42777: out <= 16'h01C9;    16'd42778: out <= 16'hFD62;    16'd42779: out <= 16'hFB37;
    16'd42780: out <= 16'hF7C6;    16'd42781: out <= 16'h05CF;    16'd42782: out <= 16'hFED1;    16'd42783: out <= 16'h01DF;
    16'd42784: out <= 16'hFFD0;    16'd42785: out <= 16'hFD77;    16'd42786: out <= 16'h00B5;    16'd42787: out <= 16'h0762;
    16'd42788: out <= 16'h0560;    16'd42789: out <= 16'h0911;    16'd42790: out <= 16'h0739;    16'd42791: out <= 16'h06FA;
    16'd42792: out <= 16'h00E4;    16'd42793: out <= 16'h0797;    16'd42794: out <= 16'hFEA2;    16'd42795: out <= 16'h0DE5;
    16'd42796: out <= 16'h0495;    16'd42797: out <= 16'h0185;    16'd42798: out <= 16'hFBF9;    16'd42799: out <= 16'h04DD;
    16'd42800: out <= 16'h0922;    16'd42801: out <= 16'h042B;    16'd42802: out <= 16'hFDCF;    16'd42803: out <= 16'h0437;
    16'd42804: out <= 16'h016C;    16'd42805: out <= 16'h08B4;    16'd42806: out <= 16'h06C2;    16'd42807: out <= 16'h0655;
    16'd42808: out <= 16'h0051;    16'd42809: out <= 16'h0539;    16'd42810: out <= 16'h0960;    16'd42811: out <= 16'h049D;
    16'd42812: out <= 16'h0149;    16'd42813: out <= 16'h03E7;    16'd42814: out <= 16'h06EE;    16'd42815: out <= 16'h06D7;
    16'd42816: out <= 16'h02C2;    16'd42817: out <= 16'h02C5;    16'd42818: out <= 16'h089D;    16'd42819: out <= 16'h0499;
    16'd42820: out <= 16'h04D8;    16'd42821: out <= 16'h0192;    16'd42822: out <= 16'hFF0A;    16'd42823: out <= 16'h07FA;
    16'd42824: out <= 16'h09BD;    16'd42825: out <= 16'hFE3F;    16'd42826: out <= 16'h0A5C;    16'd42827: out <= 16'h0350;
    16'd42828: out <= 16'h04A5;    16'd42829: out <= 16'h03F4;    16'd42830: out <= 16'hFFBF;    16'd42831: out <= 16'h0551;
    16'd42832: out <= 16'h09B7;    16'd42833: out <= 16'h03A7;    16'd42834: out <= 16'h0144;    16'd42835: out <= 16'hFEEC;
    16'd42836: out <= 16'h0520;    16'd42837: out <= 16'h01B9;    16'd42838: out <= 16'h0629;    16'd42839: out <= 16'h06CF;
    16'd42840: out <= 16'h084F;    16'd42841: out <= 16'h0322;    16'd42842: out <= 16'hFF9B;    16'd42843: out <= 16'h0033;
    16'd42844: out <= 16'hFEA5;    16'd42845: out <= 16'h057F;    16'd42846: out <= 16'h04F4;    16'd42847: out <= 16'h0639;
    16'd42848: out <= 16'h0852;    16'd42849: out <= 16'h01F3;    16'd42850: out <= 16'h076F;    16'd42851: out <= 16'h096B;
    16'd42852: out <= 16'h0626;    16'd42853: out <= 16'h02B4;    16'd42854: out <= 16'hFBC3;    16'd42855: out <= 16'h02D9;
    16'd42856: out <= 16'h03CD;    16'd42857: out <= 16'hFD1F;    16'd42858: out <= 16'h03B5;    16'd42859: out <= 16'h007E;
    16'd42860: out <= 16'h08D1;    16'd42861: out <= 16'h0041;    16'd42862: out <= 16'h03EE;    16'd42863: out <= 16'hFFEF;
    16'd42864: out <= 16'hFDD4;    16'd42865: out <= 16'hFEEF;    16'd42866: out <= 16'h050C;    16'd42867: out <= 16'h07AB;
    16'd42868: out <= 16'h02B3;    16'd42869: out <= 16'hFEDD;    16'd42870: out <= 16'h0125;    16'd42871: out <= 16'h074D;
    16'd42872: out <= 16'h07B1;    16'd42873: out <= 16'h03D8;    16'd42874: out <= 16'h095A;    16'd42875: out <= 16'h04F4;
    16'd42876: out <= 16'h0351;    16'd42877: out <= 16'hFE99;    16'd42878: out <= 16'h00E3;    16'd42879: out <= 16'hF834;
    16'd42880: out <= 16'h0385;    16'd42881: out <= 16'h0449;    16'd42882: out <= 16'h068A;    16'd42883: out <= 16'h0645;
    16'd42884: out <= 16'h01C3;    16'd42885: out <= 16'h0510;    16'd42886: out <= 16'h08A4;    16'd42887: out <= 16'h04D7;
    16'd42888: out <= 16'h01DB;    16'd42889: out <= 16'h0091;    16'd42890: out <= 16'h0740;    16'd42891: out <= 16'h05F9;
    16'd42892: out <= 16'h07D5;    16'd42893: out <= 16'h0AD9;    16'd42894: out <= 16'h053F;    16'd42895: out <= 16'h070A;
    16'd42896: out <= 16'h02F9;    16'd42897: out <= 16'hFA60;    16'd42898: out <= 16'h0459;    16'd42899: out <= 16'h0240;
    16'd42900: out <= 16'h005E;    16'd42901: out <= 16'hFF7D;    16'd42902: out <= 16'hFED8;    16'd42903: out <= 16'h06E9;
    16'd42904: out <= 16'h08BB;    16'd42905: out <= 16'h0535;    16'd42906: out <= 16'h07C0;    16'd42907: out <= 16'hFBF7;
    16'd42908: out <= 16'h03B7;    16'd42909: out <= 16'h0534;    16'd42910: out <= 16'hFDAA;    16'd42911: out <= 16'h0336;
    16'd42912: out <= 16'h05E0;    16'd42913: out <= 16'h0126;    16'd42914: out <= 16'h0541;    16'd42915: out <= 16'hFE17;
    16'd42916: out <= 16'h03C2;    16'd42917: out <= 16'h0324;    16'd42918: out <= 16'h018C;    16'd42919: out <= 16'h0095;
    16'd42920: out <= 16'h04BE;    16'd42921: out <= 16'h0516;    16'd42922: out <= 16'h01E6;    16'd42923: out <= 16'h0521;
    16'd42924: out <= 16'h0071;    16'd42925: out <= 16'hFF99;    16'd42926: out <= 16'h003C;    16'd42927: out <= 16'h07DF;
    16'd42928: out <= 16'h0564;    16'd42929: out <= 16'h05D1;    16'd42930: out <= 16'h0956;    16'd42931: out <= 16'h08AE;
    16'd42932: out <= 16'h065D;    16'd42933: out <= 16'hFF42;    16'd42934: out <= 16'h0573;    16'd42935: out <= 16'hFE0A;
    16'd42936: out <= 16'hFFA8;    16'd42937: out <= 16'hF997;    16'd42938: out <= 16'h01D1;    16'd42939: out <= 16'h059E;
    16'd42940: out <= 16'h032A;    16'd42941: out <= 16'h01CC;    16'd42942: out <= 16'hFFFF;    16'd42943: out <= 16'h00E8;
    16'd42944: out <= 16'hFCDB;    16'd42945: out <= 16'h0313;    16'd42946: out <= 16'hFE4D;    16'd42947: out <= 16'h0119;
    16'd42948: out <= 16'h039C;    16'd42949: out <= 16'hFD59;    16'd42950: out <= 16'h056B;    16'd42951: out <= 16'h05FC;
    16'd42952: out <= 16'h01F0;    16'd42953: out <= 16'h04D5;    16'd42954: out <= 16'h03B9;    16'd42955: out <= 16'h08AA;
    16'd42956: out <= 16'h0524;    16'd42957: out <= 16'h05DE;    16'd42958: out <= 16'h0670;    16'd42959: out <= 16'h05EA;
    16'd42960: out <= 16'h0318;    16'd42961: out <= 16'h080A;    16'd42962: out <= 16'h0735;    16'd42963: out <= 16'h0067;
    16'd42964: out <= 16'h037E;    16'd42965: out <= 16'h0444;    16'd42966: out <= 16'h0634;    16'd42967: out <= 16'h027E;
    16'd42968: out <= 16'h040D;    16'd42969: out <= 16'h0075;    16'd42970: out <= 16'hFA8A;    16'd42971: out <= 16'h0574;
    16'd42972: out <= 16'h046D;    16'd42973: out <= 16'hFD56;    16'd42974: out <= 16'h0400;    16'd42975: out <= 16'hFA10;
    16'd42976: out <= 16'h00B8;    16'd42977: out <= 16'hFDA3;    16'd42978: out <= 16'hFD0E;    16'd42979: out <= 16'h00E3;
    16'd42980: out <= 16'hFFD5;    16'd42981: out <= 16'h0151;    16'd42982: out <= 16'h00ED;    16'd42983: out <= 16'h0010;
    16'd42984: out <= 16'h05FD;    16'd42985: out <= 16'h004C;    16'd42986: out <= 16'h007E;    16'd42987: out <= 16'hFCBE;
    16'd42988: out <= 16'h0296;    16'd42989: out <= 16'hFCAF;    16'd42990: out <= 16'hF84D;    16'd42991: out <= 16'h00A7;
    16'd42992: out <= 16'h0444;    16'd42993: out <= 16'hFF5B;    16'd42994: out <= 16'hFE97;    16'd42995: out <= 16'h0108;
    16'd42996: out <= 16'h0166;    16'd42997: out <= 16'hFF58;    16'd42998: out <= 16'hFD73;    16'd42999: out <= 16'hF7FF;
    16'd43000: out <= 16'hF889;    16'd43001: out <= 16'h0273;    16'd43002: out <= 16'h0312;    16'd43003: out <= 16'hFC0B;
    16'd43004: out <= 16'h014D;    16'd43005: out <= 16'h0115;    16'd43006: out <= 16'hFE47;    16'd43007: out <= 16'hFC7C;
    16'd43008: out <= 16'h001C;    16'd43009: out <= 16'hFDCF;    16'd43010: out <= 16'h00E5;    16'd43011: out <= 16'h0212;
    16'd43012: out <= 16'h0279;    16'd43013: out <= 16'hFEE6;    16'd43014: out <= 16'h005B;    16'd43015: out <= 16'h02A0;
    16'd43016: out <= 16'h05C9;    16'd43017: out <= 16'hFDBE;    16'd43018: out <= 16'hFD28;    16'd43019: out <= 16'hF7A9;
    16'd43020: out <= 16'h043B;    16'd43021: out <= 16'h0046;    16'd43022: out <= 16'h04DA;    16'd43023: out <= 16'h042D;
    16'd43024: out <= 16'hF7E3;    16'd43025: out <= 16'h02DA;    16'd43026: out <= 16'h002F;    16'd43027: out <= 16'h00F2;
    16'd43028: out <= 16'h029D;    16'd43029: out <= 16'h00C6;    16'd43030: out <= 16'hFFE2;    16'd43031: out <= 16'h01BB;
    16'd43032: out <= 16'h0014;    16'd43033: out <= 16'h0291;    16'd43034: out <= 16'hF9DB;    16'd43035: out <= 16'h029C;
    16'd43036: out <= 16'h0077;    16'd43037: out <= 16'hFA9B;    16'd43038: out <= 16'hFDCA;    16'd43039: out <= 16'hFCF9;
    16'd43040: out <= 16'h04EB;    16'd43041: out <= 16'h0339;    16'd43042: out <= 16'h01BC;    16'd43043: out <= 16'h0552;
    16'd43044: out <= 16'h0588;    16'd43045: out <= 16'hFF73;    16'd43046: out <= 16'h095C;    16'd43047: out <= 16'h06DE;
    16'd43048: out <= 16'h03C6;    16'd43049: out <= 16'h07A6;    16'd43050: out <= 16'h013D;    16'd43051: out <= 16'h041A;
    16'd43052: out <= 16'h02F7;    16'd43053: out <= 16'h06DF;    16'd43054: out <= 16'h09E8;    16'd43055: out <= 16'h0CAD;
    16'd43056: out <= 16'hFEBD;    16'd43057: out <= 16'h0607;    16'd43058: out <= 16'hFAF6;    16'd43059: out <= 16'h03B0;
    16'd43060: out <= 16'h01DB;    16'd43061: out <= 16'h026D;    16'd43062: out <= 16'h0476;    16'd43063: out <= 16'h0848;
    16'd43064: out <= 16'h0182;    16'd43065: out <= 16'h0401;    16'd43066: out <= 16'h03CD;    16'd43067: out <= 16'hFE0D;
    16'd43068: out <= 16'h02EA;    16'd43069: out <= 16'h0054;    16'd43070: out <= 16'h0309;    16'd43071: out <= 16'hFF6B;
    16'd43072: out <= 16'h0846;    16'd43073: out <= 16'h0975;    16'd43074: out <= 16'hFF3C;    16'd43075: out <= 16'h0045;
    16'd43076: out <= 16'h0805;    16'd43077: out <= 16'h0022;    16'd43078: out <= 16'hFDF2;    16'd43079: out <= 16'h0036;
    16'd43080: out <= 16'h0118;    16'd43081: out <= 16'h0363;    16'd43082: out <= 16'hFB6A;    16'd43083: out <= 16'h0609;
    16'd43084: out <= 16'h080B;    16'd43085: out <= 16'h0555;    16'd43086: out <= 16'h08B3;    16'd43087: out <= 16'h00A2;
    16'd43088: out <= 16'h0AE3;    16'd43089: out <= 16'h07BC;    16'd43090: out <= 16'h0884;    16'd43091: out <= 16'h051E;
    16'd43092: out <= 16'h0AE8;    16'd43093: out <= 16'h010F;    16'd43094: out <= 16'h0833;    16'd43095: out <= 16'h0215;
    16'd43096: out <= 16'hF8A1;    16'd43097: out <= 16'h056C;    16'd43098: out <= 16'h0341;    16'd43099: out <= 16'h072D;
    16'd43100: out <= 16'hFFFD;    16'd43101: out <= 16'hFE8F;    16'd43102: out <= 16'h0302;    16'd43103: out <= 16'h0962;
    16'd43104: out <= 16'h01C9;    16'd43105: out <= 16'h0589;    16'd43106: out <= 16'h06E2;    16'd43107: out <= 16'h08E5;
    16'd43108: out <= 16'h034B;    16'd43109: out <= 16'hFE42;    16'd43110: out <= 16'h0450;    16'd43111: out <= 16'h0C2E;
    16'd43112: out <= 16'h0243;    16'd43113: out <= 16'h04C2;    16'd43114: out <= 16'h0100;    16'd43115: out <= 16'hFBFA;
    16'd43116: out <= 16'h06AA;    16'd43117: out <= 16'h019B;    16'd43118: out <= 16'h0706;    16'd43119: out <= 16'h0BEC;
    16'd43120: out <= 16'h0C86;    16'd43121: out <= 16'h03CC;    16'd43122: out <= 16'hF871;    16'd43123: out <= 16'h0743;
    16'd43124: out <= 16'h016B;    16'd43125: out <= 16'h09BE;    16'd43126: out <= 16'h045C;    16'd43127: out <= 16'h0467;
    16'd43128: out <= 16'hFF5F;    16'd43129: out <= 16'h0BDC;    16'd43130: out <= 16'h0143;    16'd43131: out <= 16'h0558;
    16'd43132: out <= 16'hFE64;    16'd43133: out <= 16'h0A30;    16'd43134: out <= 16'h03B3;    16'd43135: out <= 16'h0472;
    16'd43136: out <= 16'h0379;    16'd43137: out <= 16'hFE0D;    16'd43138: out <= 16'h05F7;    16'd43139: out <= 16'h0413;
    16'd43140: out <= 16'h0306;    16'd43141: out <= 16'h0A72;    16'd43142: out <= 16'h009B;    16'd43143: out <= 16'h0010;
    16'd43144: out <= 16'h01B5;    16'd43145: out <= 16'h03D1;    16'd43146: out <= 16'h0BCD;    16'd43147: out <= 16'h0076;
    16'd43148: out <= 16'h04A8;    16'd43149: out <= 16'h0607;    16'd43150: out <= 16'h04B2;    16'd43151: out <= 16'h017A;
    16'd43152: out <= 16'hFE97;    16'd43153: out <= 16'h0260;    16'd43154: out <= 16'h088B;    16'd43155: out <= 16'h0108;
    16'd43156: out <= 16'h0975;    16'd43157: out <= 16'h0743;    16'd43158: out <= 16'h0814;    16'd43159: out <= 16'h0123;
    16'd43160: out <= 16'h0547;    16'd43161: out <= 16'h0242;    16'd43162: out <= 16'h0700;    16'd43163: out <= 16'h06D2;
    16'd43164: out <= 16'h0118;    16'd43165: out <= 16'hFDF7;    16'd43166: out <= 16'hFFC0;    16'd43167: out <= 16'h079E;
    16'd43168: out <= 16'h0BB8;    16'd43169: out <= 16'h033E;    16'd43170: out <= 16'hFF81;    16'd43171: out <= 16'hF7F7;
    16'd43172: out <= 16'h05A8;    16'd43173: out <= 16'h048B;    16'd43174: out <= 16'h0508;    16'd43175: out <= 16'h0620;
    16'd43176: out <= 16'h091C;    16'd43177: out <= 16'h065D;    16'd43178: out <= 16'h0761;    16'd43179: out <= 16'h0232;
    16'd43180: out <= 16'hFC28;    16'd43181: out <= 16'h0714;    16'd43182: out <= 16'h06FB;    16'd43183: out <= 16'h0375;
    16'd43184: out <= 16'h0385;    16'd43185: out <= 16'h0234;    16'd43186: out <= 16'h0B61;    16'd43187: out <= 16'h0AE9;
    16'd43188: out <= 16'h0153;    16'd43189: out <= 16'hFDB5;    16'd43190: out <= 16'h0482;    16'd43191: out <= 16'h06F1;
    16'd43192: out <= 16'h02B1;    16'd43193: out <= 16'h05B4;    16'd43194: out <= 16'h082F;    16'd43195: out <= 16'hFD1C;
    16'd43196: out <= 16'hFCEF;    16'd43197: out <= 16'h0968;    16'd43198: out <= 16'h00C9;    16'd43199: out <= 16'h069B;
    16'd43200: out <= 16'h03B7;    16'd43201: out <= 16'h0729;    16'd43202: out <= 16'h0428;    16'd43203: out <= 16'h0A39;
    16'd43204: out <= 16'h048A;    16'd43205: out <= 16'h09A6;    16'd43206: out <= 16'h070F;    16'd43207: out <= 16'h03FB;
    16'd43208: out <= 16'h0D0F;    16'd43209: out <= 16'hFDBB;    16'd43210: out <= 16'h0714;    16'd43211: out <= 16'h04FC;
    16'd43212: out <= 16'h0263;    16'd43213: out <= 16'hFED4;    16'd43214: out <= 16'h0108;    16'd43215: out <= 16'h024B;
    16'd43216: out <= 16'h0153;    16'd43217: out <= 16'h0054;    16'd43218: out <= 16'hFF96;    16'd43219: out <= 16'h03E7;
    16'd43220: out <= 16'h0567;    16'd43221: out <= 16'hFF8F;    16'd43222: out <= 16'h0372;    16'd43223: out <= 16'h040F;
    16'd43224: out <= 16'h0273;    16'd43225: out <= 16'h01E3;    16'd43226: out <= 16'h0935;    16'd43227: out <= 16'hF87D;
    16'd43228: out <= 16'hFF35;    16'd43229: out <= 16'hFE6F;    16'd43230: out <= 16'hFFB8;    16'd43231: out <= 16'h001E;
    16'd43232: out <= 16'h02F4;    16'd43233: out <= 16'hFF10;    16'd43234: out <= 16'h0442;    16'd43235: out <= 16'hFE7D;
    16'd43236: out <= 16'h051A;    16'd43237: out <= 16'h00A0;    16'd43238: out <= 16'hFFAF;    16'd43239: out <= 16'h0194;
    16'd43240: out <= 16'hFC5F;    16'd43241: out <= 16'hFBDC;    16'd43242: out <= 16'hFF9B;    16'd43243: out <= 16'hFFDB;
    16'd43244: out <= 16'hFDD8;    16'd43245: out <= 16'h002F;    16'd43246: out <= 16'h0051;    16'd43247: out <= 16'hFCC3;
    16'd43248: out <= 16'hF21D;    16'd43249: out <= 16'h0138;    16'd43250: out <= 16'hFD78;    16'd43251: out <= 16'h0050;
    16'd43252: out <= 16'hF625;    16'd43253: out <= 16'h033F;    16'd43254: out <= 16'hFEED;    16'd43255: out <= 16'hFF0C;
    16'd43256: out <= 16'hFDF4;    16'd43257: out <= 16'h0168;    16'd43258: out <= 16'hFE9F;    16'd43259: out <= 16'h00EF;
    16'd43260: out <= 16'h03EB;    16'd43261: out <= 16'h0404;    16'd43262: out <= 16'h01DF;    16'd43263: out <= 16'hFD92;
    16'd43264: out <= 16'hFC31;    16'd43265: out <= 16'h0164;    16'd43266: out <= 16'h01E9;    16'd43267: out <= 16'h04A7;
    16'd43268: out <= 16'hFA1A;    16'd43269: out <= 16'hFDCA;    16'd43270: out <= 16'hFFB9;    16'd43271: out <= 16'h040D;
    16'd43272: out <= 16'h00D5;    16'd43273: out <= 16'h004C;    16'd43274: out <= 16'hFED9;    16'd43275: out <= 16'hFC66;
    16'd43276: out <= 16'h0186;    16'd43277: out <= 16'hFC9C;    16'd43278: out <= 16'hFECC;    16'd43279: out <= 16'h0176;
    16'd43280: out <= 16'hFF75;    16'd43281: out <= 16'hFE24;    16'd43282: out <= 16'hFC7A;    16'd43283: out <= 16'h0344;
    16'd43284: out <= 16'h0395;    16'd43285: out <= 16'h004E;    16'd43286: out <= 16'hFFE9;    16'd43287: out <= 16'h0501;
    16'd43288: out <= 16'h02F4;    16'd43289: out <= 16'h003A;    16'd43290: out <= 16'h00A1;    16'd43291: out <= 16'h047B;
    16'd43292: out <= 16'h0203;    16'd43293: out <= 16'hFD38;    16'd43294: out <= 16'hFEB6;    16'd43295: out <= 16'hF6FA;
    16'd43296: out <= 16'h0555;    16'd43297: out <= 16'hFFB6;    16'd43298: out <= 16'h05E8;    16'd43299: out <= 16'h06C2;
    16'd43300: out <= 16'h0617;    16'd43301: out <= 16'h0154;    16'd43302: out <= 16'h03CC;    16'd43303: out <= 16'h04F9;
    16'd43304: out <= 16'hF8F3;    16'd43305: out <= 16'h0864;    16'd43306: out <= 16'h0039;    16'd43307: out <= 16'h06C6;
    16'd43308: out <= 16'h040A;    16'd43309: out <= 16'h002E;    16'd43310: out <= 16'hFF4D;    16'd43311: out <= 16'h0435;
    16'd43312: out <= 16'h06E4;    16'd43313: out <= 16'h08CB;    16'd43314: out <= 16'h0051;    16'd43315: out <= 16'h01F3;
    16'd43316: out <= 16'hFF57;    16'd43317: out <= 16'h0562;    16'd43318: out <= 16'h0160;    16'd43319: out <= 16'h0545;
    16'd43320: out <= 16'h06DB;    16'd43321: out <= 16'h0049;    16'd43322: out <= 16'h0223;    16'd43323: out <= 16'h0287;
    16'd43324: out <= 16'hFF8C;    16'd43325: out <= 16'h017A;    16'd43326: out <= 16'h06AF;    16'd43327: out <= 16'hFF01;
    16'd43328: out <= 16'h03B9;    16'd43329: out <= 16'hFF34;    16'd43330: out <= 16'h0611;    16'd43331: out <= 16'hFB8B;
    16'd43332: out <= 16'h0526;    16'd43333: out <= 16'h017D;    16'd43334: out <= 16'h0004;    16'd43335: out <= 16'h0004;
    16'd43336: out <= 16'h0744;    16'd43337: out <= 16'h07C1;    16'd43338: out <= 16'h04C5;    16'd43339: out <= 16'h0663;
    16'd43340: out <= 16'h0527;    16'd43341: out <= 16'hFBCB;    16'd43342: out <= 16'h0471;    16'd43343: out <= 16'h015A;
    16'd43344: out <= 16'h0548;    16'd43345: out <= 16'h0393;    16'd43346: out <= 16'hFFB3;    16'd43347: out <= 16'h092A;
    16'd43348: out <= 16'hFF46;    16'd43349: out <= 16'h05C9;    16'd43350: out <= 16'h025E;    16'd43351: out <= 16'h0AFE;
    16'd43352: out <= 16'h02E8;    16'd43353: out <= 16'h0212;    16'd43354: out <= 16'h07F5;    16'd43355: out <= 16'h0B91;
    16'd43356: out <= 16'h042C;    16'd43357: out <= 16'hFB43;    16'd43358: out <= 16'h0473;    16'd43359: out <= 16'h055E;
    16'd43360: out <= 16'hFF60;    16'd43361: out <= 16'h03BB;    16'd43362: out <= 16'h01F6;    16'd43363: out <= 16'hFD34;
    16'd43364: out <= 16'h0447;    16'd43365: out <= 16'h00C6;    16'd43366: out <= 16'h031F;    16'd43367: out <= 16'hFF11;
    16'd43368: out <= 16'hFDA3;    16'd43369: out <= 16'h0603;    16'd43370: out <= 16'hFD7B;    16'd43371: out <= 16'h038A;
    16'd43372: out <= 16'h0D77;    16'd43373: out <= 16'h077C;    16'd43374: out <= 16'h0821;    16'd43375: out <= 16'h05E3;
    16'd43376: out <= 16'hFEDC;    16'd43377: out <= 16'hFD15;    16'd43378: out <= 16'h06AD;    16'd43379: out <= 16'hFDA6;
    16'd43380: out <= 16'h03D2;    16'd43381: out <= 16'h0185;    16'd43382: out <= 16'hFE30;    16'd43383: out <= 16'h054C;
    16'd43384: out <= 16'h0235;    16'd43385: out <= 16'h086C;    16'd43386: out <= 16'h0917;    16'd43387: out <= 16'h0617;
    16'd43388: out <= 16'h01F7;    16'd43389: out <= 16'h0507;    16'd43390: out <= 16'hFDC7;    16'd43391: out <= 16'h0792;
    16'd43392: out <= 16'hFED1;    16'd43393: out <= 16'h01E3;    16'd43394: out <= 16'h052E;    16'd43395: out <= 16'h0390;
    16'd43396: out <= 16'h0616;    16'd43397: out <= 16'h0CD7;    16'd43398: out <= 16'h07F7;    16'd43399: out <= 16'hFFBB;
    16'd43400: out <= 16'h084A;    16'd43401: out <= 16'h015E;    16'd43402: out <= 16'h03E0;    16'd43403: out <= 16'h0469;
    16'd43404: out <= 16'hFEC1;    16'd43405: out <= 16'h0490;    16'd43406: out <= 16'h0803;    16'd43407: out <= 16'h0367;
    16'd43408: out <= 16'h075F;    16'd43409: out <= 16'h0275;    16'd43410: out <= 16'h0903;    16'd43411: out <= 16'hFE1B;
    16'd43412: out <= 16'h05E4;    16'd43413: out <= 16'h067B;    16'd43414: out <= 16'h08F6;    16'd43415: out <= 16'h0EDB;
    16'd43416: out <= 16'hF8B4;    16'd43417: out <= 16'h02D5;    16'd43418: out <= 16'h0500;    16'd43419: out <= 16'h092E;
    16'd43420: out <= 16'h0AA9;    16'd43421: out <= 16'h02B1;    16'd43422: out <= 16'h0265;    16'd43423: out <= 16'h05EF;
    16'd43424: out <= 16'h0709;    16'd43425: out <= 16'h0C55;    16'd43426: out <= 16'hFEC8;    16'd43427: out <= 16'h0784;
    16'd43428: out <= 16'h0931;    16'd43429: out <= 16'h00C1;    16'd43430: out <= 16'h01D7;    16'd43431: out <= 16'h0798;
    16'd43432: out <= 16'h0196;    16'd43433: out <= 16'h01B4;    16'd43434: out <= 16'h0589;    16'd43435: out <= 16'h04FA;
    16'd43436: out <= 16'h04FD;    16'd43437: out <= 16'h0187;    16'd43438: out <= 16'h0162;    16'd43439: out <= 16'hFE7D;
    16'd43440: out <= 16'h0029;    16'd43441: out <= 16'h0487;    16'd43442: out <= 16'h0223;    16'd43443: out <= 16'h01B3;
    16'd43444: out <= 16'h00E5;    16'd43445: out <= 16'h0C73;    16'd43446: out <= 16'h05EF;    16'd43447: out <= 16'hFC86;
    16'd43448: out <= 16'h04F1;    16'd43449: out <= 16'hFC58;    16'd43450: out <= 16'h0043;    16'd43451: out <= 16'h02F7;
    16'd43452: out <= 16'h06FA;    16'd43453: out <= 16'h0AEA;    16'd43454: out <= 16'hFD84;    16'd43455: out <= 16'h0515;
    16'd43456: out <= 16'h0451;    16'd43457: out <= 16'h09D9;    16'd43458: out <= 16'h0153;    16'd43459: out <= 16'h033A;
    16'd43460: out <= 16'h040B;    16'd43461: out <= 16'h02D6;    16'd43462: out <= 16'h09B4;    16'd43463: out <= 16'hF86D;
    16'd43464: out <= 16'h033D;    16'd43465: out <= 16'hFF7C;    16'd43466: out <= 16'hFE75;    16'd43467: out <= 16'h06B3;
    16'd43468: out <= 16'h0496;    16'd43469: out <= 16'h06BB;    16'd43470: out <= 16'h06D9;    16'd43471: out <= 16'h0971;
    16'd43472: out <= 16'h033E;    16'd43473: out <= 16'h0122;    16'd43474: out <= 16'h045A;    16'd43475: out <= 16'h06D7;
    16'd43476: out <= 16'h05DD;    16'd43477: out <= 16'h04FC;    16'd43478: out <= 16'hFDC3;    16'd43479: out <= 16'hFF65;
    16'd43480: out <= 16'h01CC;    16'd43481: out <= 16'h0257;    16'd43482: out <= 16'h059E;    16'd43483: out <= 16'hFCEC;
    16'd43484: out <= 16'hFD02;    16'd43485: out <= 16'hFB62;    16'd43486: out <= 16'hF9E5;    16'd43487: out <= 16'h006A;
    16'd43488: out <= 16'hFEE6;    16'd43489: out <= 16'h0129;    16'd43490: out <= 16'h03C5;    16'd43491: out <= 16'h0172;
    16'd43492: out <= 16'hFBBC;    16'd43493: out <= 16'h02B8;    16'd43494: out <= 16'hFB22;    16'd43495: out <= 16'hFEEA;
    16'd43496: out <= 16'h04BB;    16'd43497: out <= 16'h0179;    16'd43498: out <= 16'h0321;    16'd43499: out <= 16'h05D7;
    16'd43500: out <= 16'h02EE;    16'd43501: out <= 16'h0071;    16'd43502: out <= 16'h0740;    16'd43503: out <= 16'hFDA7;
    16'd43504: out <= 16'h03E1;    16'd43505: out <= 16'h0080;    16'd43506: out <= 16'hFEC1;    16'd43507: out <= 16'h019F;
    16'd43508: out <= 16'h0352;    16'd43509: out <= 16'hFD11;    16'd43510: out <= 16'hFFB8;    16'd43511: out <= 16'h01C4;
    16'd43512: out <= 16'h0301;    16'd43513: out <= 16'hFACB;    16'd43514: out <= 16'hFDA5;    16'd43515: out <= 16'hFFC4;
    16'd43516: out <= 16'h0246;    16'd43517: out <= 16'hFE25;    16'd43518: out <= 16'hFECB;    16'd43519: out <= 16'hFBE6;
    16'd43520: out <= 16'h06FD;    16'd43521: out <= 16'h0224;    16'd43522: out <= 16'h013C;    16'd43523: out <= 16'h0410;
    16'd43524: out <= 16'h04FF;    16'd43525: out <= 16'h04F3;    16'd43526: out <= 16'h0471;    16'd43527: out <= 16'hFE7E;
    16'd43528: out <= 16'h01B3;    16'd43529: out <= 16'hFE2E;    16'd43530: out <= 16'h0117;    16'd43531: out <= 16'h0475;
    16'd43532: out <= 16'hFEF6;    16'd43533: out <= 16'hFD24;    16'd43534: out <= 16'h00CA;    16'd43535: out <= 16'hFBE1;
    16'd43536: out <= 16'hFD3B;    16'd43537: out <= 16'hFEB3;    16'd43538: out <= 16'hFEB2;    16'd43539: out <= 16'hFDC2;
    16'd43540: out <= 16'h06AB;    16'd43541: out <= 16'h08AE;    16'd43542: out <= 16'h040B;    16'd43543: out <= 16'h0550;
    16'd43544: out <= 16'h02C5;    16'd43545: out <= 16'hFF99;    16'd43546: out <= 16'hFCEA;    16'd43547: out <= 16'h06E6;
    16'd43548: out <= 16'hFF59;    16'd43549: out <= 16'hFACD;    16'd43550: out <= 16'hFF02;    16'd43551: out <= 16'h00AE;
    16'd43552: out <= 16'hFC51;    16'd43553: out <= 16'h012E;    16'd43554: out <= 16'h0708;    16'd43555: out <= 16'h01B6;
    16'd43556: out <= 16'h03FF;    16'd43557: out <= 16'h0101;    16'd43558: out <= 16'h0C6A;    16'd43559: out <= 16'h0533;
    16'd43560: out <= 16'hFE3F;    16'd43561: out <= 16'h01C6;    16'd43562: out <= 16'hF8BF;    16'd43563: out <= 16'h03D4;
    16'd43564: out <= 16'h03A7;    16'd43565: out <= 16'h0333;    16'd43566: out <= 16'h0381;    16'd43567: out <= 16'h087B;
    16'd43568: out <= 16'h0527;    16'd43569: out <= 16'h089B;    16'd43570: out <= 16'hFA24;    16'd43571: out <= 16'h0AE1;
    16'd43572: out <= 16'h132F;    16'd43573: out <= 16'h064B;    16'd43574: out <= 16'hFA47;    16'd43575: out <= 16'h060C;
    16'd43576: out <= 16'h0502;    16'd43577: out <= 16'h05AA;    16'd43578: out <= 16'h0461;    16'd43579: out <= 16'h05F2;
    16'd43580: out <= 16'hF9ED;    16'd43581: out <= 16'h097D;    16'd43582: out <= 16'h0D4A;    16'd43583: out <= 16'h0203;
    16'd43584: out <= 16'hFAB4;    16'd43585: out <= 16'h02A9;    16'd43586: out <= 16'h0827;    16'd43587: out <= 16'h00E2;
    16'd43588: out <= 16'h0387;    16'd43589: out <= 16'h0A13;    16'd43590: out <= 16'h0417;    16'd43591: out <= 16'h0468;
    16'd43592: out <= 16'h0C75;    16'd43593: out <= 16'h01C0;    16'd43594: out <= 16'hFF7D;    16'd43595: out <= 16'h029F;
    16'd43596: out <= 16'h08BB;    16'd43597: out <= 16'h0354;    16'd43598: out <= 16'h02BE;    16'd43599: out <= 16'h05DC;
    16'd43600: out <= 16'h019B;    16'd43601: out <= 16'h06BF;    16'd43602: out <= 16'h08F8;    16'd43603: out <= 16'h03B6;
    16'd43604: out <= 16'h03A7;    16'd43605: out <= 16'h058D;    16'd43606: out <= 16'h03AC;    16'd43607: out <= 16'h0483;
    16'd43608: out <= 16'h04B0;    16'd43609: out <= 16'h0366;    16'd43610: out <= 16'h03FF;    16'd43611: out <= 16'h04DB;
    16'd43612: out <= 16'h01A1;    16'd43613: out <= 16'h06F8;    16'd43614: out <= 16'h0017;    16'd43615: out <= 16'h085E;
    16'd43616: out <= 16'h08C3;    16'd43617: out <= 16'h0402;    16'd43618: out <= 16'h0647;    16'd43619: out <= 16'h0401;
    16'd43620: out <= 16'h064A;    16'd43621: out <= 16'h03CA;    16'd43622: out <= 16'h02E3;    16'd43623: out <= 16'h06BD;
    16'd43624: out <= 16'h07F7;    16'd43625: out <= 16'h082B;    16'd43626: out <= 16'h015F;    16'd43627: out <= 16'h089D;
    16'd43628: out <= 16'hFF95;    16'd43629: out <= 16'h02C1;    16'd43630: out <= 16'h06CC;    16'd43631: out <= 16'h0079;
    16'd43632: out <= 16'h0077;    16'd43633: out <= 16'h070F;    16'd43634: out <= 16'hFC3D;    16'd43635: out <= 16'hFFC5;
    16'd43636: out <= 16'h0261;    16'd43637: out <= 16'h0D0D;    16'd43638: out <= 16'h041B;    16'd43639: out <= 16'h0502;
    16'd43640: out <= 16'h06D4;    16'd43641: out <= 16'h0741;    16'd43642: out <= 16'h06AD;    16'd43643: out <= 16'h058F;
    16'd43644: out <= 16'h02EC;    16'd43645: out <= 16'h09C5;    16'd43646: out <= 16'hFFD6;    16'd43647: out <= 16'h022D;
    16'd43648: out <= 16'hFF9F;    16'd43649: out <= 16'hFBFD;    16'd43650: out <= 16'h0C56;    16'd43651: out <= 16'h0251;
    16'd43652: out <= 16'h044D;    16'd43653: out <= 16'h05A9;    16'd43654: out <= 16'h0714;    16'd43655: out <= 16'h03D4;
    16'd43656: out <= 16'h0133;    16'd43657: out <= 16'h0089;    16'd43658: out <= 16'h0335;    16'd43659: out <= 16'h044E;
    16'd43660: out <= 16'h0009;    16'd43661: out <= 16'h064D;    16'd43662: out <= 16'h07C3;    16'd43663: out <= 16'h05CD;
    16'd43664: out <= 16'h04BE;    16'd43665: out <= 16'h0146;    16'd43666: out <= 16'h02B8;    16'd43667: out <= 16'h01F3;
    16'd43668: out <= 16'h0117;    16'd43669: out <= 16'h0B3B;    16'd43670: out <= 16'h00D3;    16'd43671: out <= 16'hFE38;
    16'd43672: out <= 16'h07AD;    16'd43673: out <= 16'h0329;    16'd43674: out <= 16'hFFDB;    16'd43675: out <= 16'h0933;
    16'd43676: out <= 16'h0351;    16'd43677: out <= 16'h069D;    16'd43678: out <= 16'h0453;    16'd43679: out <= 16'h0952;
    16'd43680: out <= 16'h08C5;    16'd43681: out <= 16'h08D9;    16'd43682: out <= 16'h0634;    16'd43683: out <= 16'h050A;
    16'd43684: out <= 16'h016E;    16'd43685: out <= 16'h0557;    16'd43686: out <= 16'h04DD;    16'd43687: out <= 16'h0036;
    16'd43688: out <= 16'h049C;    16'd43689: out <= 16'h04F9;    16'd43690: out <= 16'h043D;    16'd43691: out <= 16'h0073;
    16'd43692: out <= 16'h04E2;    16'd43693: out <= 16'h00AF;    16'd43694: out <= 16'h0832;    16'd43695: out <= 16'h0402;
    16'd43696: out <= 16'h0511;    16'd43697: out <= 16'h061F;    16'd43698: out <= 16'h02DF;    16'd43699: out <= 16'h0902;
    16'd43700: out <= 16'h094E;    16'd43701: out <= 16'h031A;    16'd43702: out <= 16'h0597;    16'd43703: out <= 16'h026E;
    16'd43704: out <= 16'hFF71;    16'd43705: out <= 16'h0830;    16'd43706: out <= 16'hFE5F;    16'd43707: out <= 16'h0166;
    16'd43708: out <= 16'h03C2;    16'd43709: out <= 16'h083F;    16'd43710: out <= 16'hFE2C;    16'd43711: out <= 16'h03B5;
    16'd43712: out <= 16'h0117;    16'd43713: out <= 16'h03C8;    16'd43714: out <= 16'h00C5;    16'd43715: out <= 16'h0470;
    16'd43716: out <= 16'hFFE6;    16'd43717: out <= 16'h023D;    16'd43718: out <= 16'h0583;    16'd43719: out <= 16'hFDFA;
    16'd43720: out <= 16'h045E;    16'd43721: out <= 16'h0AA6;    16'd43722: out <= 16'h055D;    16'd43723: out <= 16'h029E;
    16'd43724: out <= 16'h07D1;    16'd43725: out <= 16'h0A00;    16'd43726: out <= 16'h02E9;    16'd43727: out <= 16'h0344;
    16'd43728: out <= 16'h00F8;    16'd43729: out <= 16'h0634;    16'd43730: out <= 16'h069B;    16'd43731: out <= 16'h02AC;
    16'd43732: out <= 16'h0865;    16'd43733: out <= 16'h05AE;    16'd43734: out <= 16'hFB5A;    16'd43735: out <= 16'hFBA7;
    16'd43736: out <= 16'h03DD;    16'd43737: out <= 16'h00BD;    16'd43738: out <= 16'hFDEB;    16'd43739: out <= 16'hFE6E;
    16'd43740: out <= 16'h014F;    16'd43741: out <= 16'h048F;    16'd43742: out <= 16'h02B3;    16'd43743: out <= 16'h012C;
    16'd43744: out <= 16'h01EE;    16'd43745: out <= 16'hFDFE;    16'd43746: out <= 16'h068C;    16'd43747: out <= 16'h02E9;
    16'd43748: out <= 16'hFCA6;    16'd43749: out <= 16'h0405;    16'd43750: out <= 16'h060C;    16'd43751: out <= 16'h036C;
    16'd43752: out <= 16'hFE0B;    16'd43753: out <= 16'hFD24;    16'd43754: out <= 16'h01CA;    16'd43755: out <= 16'h021E;
    16'd43756: out <= 16'hFF0B;    16'd43757: out <= 16'h071E;    16'd43758: out <= 16'hFF91;    16'd43759: out <= 16'h00F4;
    16'd43760: out <= 16'h0336;    16'd43761: out <= 16'h0200;    16'd43762: out <= 16'h0260;    16'd43763: out <= 16'h0966;
    16'd43764: out <= 16'h0021;    16'd43765: out <= 16'h0290;    16'd43766: out <= 16'hFFA3;    16'd43767: out <= 16'hFDC8;
    16'd43768: out <= 16'h011C;    16'd43769: out <= 16'h0110;    16'd43770: out <= 16'h015E;    16'd43771: out <= 16'h014B;
    16'd43772: out <= 16'h01CC;    16'd43773: out <= 16'hFEC7;    16'd43774: out <= 16'hFD60;    16'd43775: out <= 16'h023B;
    16'd43776: out <= 16'hFF68;    16'd43777: out <= 16'hF9CF;    16'd43778: out <= 16'hFC4D;    16'd43779: out <= 16'hFC14;
    16'd43780: out <= 16'hFDDC;    16'd43781: out <= 16'hFF66;    16'd43782: out <= 16'h0111;    16'd43783: out <= 16'hFFE7;
    16'd43784: out <= 16'hFCCC;    16'd43785: out <= 16'h0602;    16'd43786: out <= 16'hFDC9;    16'd43787: out <= 16'hFF4D;
    16'd43788: out <= 16'h0336;    16'd43789: out <= 16'hFBA3;    16'd43790: out <= 16'hFECE;    16'd43791: out <= 16'h00CF;
    16'd43792: out <= 16'h065A;    16'd43793: out <= 16'hFD9B;    16'd43794: out <= 16'hFCFC;    16'd43795: out <= 16'hFD01;
    16'd43796: out <= 16'hFD0A;    16'd43797: out <= 16'h0016;    16'd43798: out <= 16'h04DA;    16'd43799: out <= 16'hFADF;
    16'd43800: out <= 16'h0A20;    16'd43801: out <= 16'hF890;    16'd43802: out <= 16'h003D;    16'd43803: out <= 16'hFDE2;
    16'd43804: out <= 16'h04D7;    16'd43805: out <= 16'hFA8E;    16'd43806: out <= 16'hFF18;    16'd43807: out <= 16'h068A;
    16'd43808: out <= 16'hFCF0;    16'd43809: out <= 16'h0040;    16'd43810: out <= 16'h068A;    16'd43811: out <= 16'hFE1D;
    16'd43812: out <= 16'h015A;    16'd43813: out <= 16'h08AC;    16'd43814: out <= 16'h04AB;    16'd43815: out <= 16'h0965;
    16'd43816: out <= 16'h0719;    16'd43817: out <= 16'h0113;    16'd43818: out <= 16'hFFA8;    16'd43819: out <= 16'h079A;
    16'd43820: out <= 16'h031A;    16'd43821: out <= 16'h0514;    16'd43822: out <= 16'h02E1;    16'd43823: out <= 16'h0575;
    16'd43824: out <= 16'h036F;    16'd43825: out <= 16'h0274;    16'd43826: out <= 16'h0B67;    16'd43827: out <= 16'h043D;
    16'd43828: out <= 16'h09FC;    16'd43829: out <= 16'h00A3;    16'd43830: out <= 16'h0783;    16'd43831: out <= 16'h02F2;
    16'd43832: out <= 16'h03A2;    16'd43833: out <= 16'h01D3;    16'd43834: out <= 16'h06CE;    16'd43835: out <= 16'h00B0;
    16'd43836: out <= 16'h0A8E;    16'd43837: out <= 16'h0614;    16'd43838: out <= 16'hFC48;    16'd43839: out <= 16'h0AFD;
    16'd43840: out <= 16'h03F0;    16'd43841: out <= 16'h015D;    16'd43842: out <= 16'hFF58;    16'd43843: out <= 16'h0821;
    16'd43844: out <= 16'h0335;    16'd43845: out <= 16'h047B;    16'd43846: out <= 16'hFFAB;    16'd43847: out <= 16'h03B2;
    16'd43848: out <= 16'h0DEA;    16'd43849: out <= 16'hFE02;    16'd43850: out <= 16'h0249;    16'd43851: out <= 16'h031F;
    16'd43852: out <= 16'h09AF;    16'd43853: out <= 16'h006D;    16'd43854: out <= 16'hFF4E;    16'd43855: out <= 16'hFE4D;
    16'd43856: out <= 16'h03BD;    16'd43857: out <= 16'h0265;    16'd43858: out <= 16'h02C2;    16'd43859: out <= 16'h0529;
    16'd43860: out <= 16'h0205;    16'd43861: out <= 16'h0455;    16'd43862: out <= 16'h04E0;    16'd43863: out <= 16'h024C;
    16'd43864: out <= 16'h034E;    16'd43865: out <= 16'h01D8;    16'd43866: out <= 16'h0287;    16'd43867: out <= 16'h0117;
    16'd43868: out <= 16'h096E;    16'd43869: out <= 16'h04FA;    16'd43870: out <= 16'h0258;    16'd43871: out <= 16'h051B;
    16'd43872: out <= 16'h08E2;    16'd43873: out <= 16'hFFE9;    16'd43874: out <= 16'h05E3;    16'd43875: out <= 16'h0821;
    16'd43876: out <= 16'h01B6;    16'd43877: out <= 16'h0433;    16'd43878: out <= 16'h0BA0;    16'd43879: out <= 16'h01E2;
    16'd43880: out <= 16'h008B;    16'd43881: out <= 16'h048B;    16'd43882: out <= 16'hFC20;    16'd43883: out <= 16'h076C;
    16'd43884: out <= 16'h00A5;    16'd43885: out <= 16'h0AB3;    16'd43886: out <= 16'h06E7;    16'd43887: out <= 16'h0473;
    16'd43888: out <= 16'h01BA;    16'd43889: out <= 16'h0625;    16'd43890: out <= 16'h0475;    16'd43891: out <= 16'h0740;
    16'd43892: out <= 16'h0083;    16'd43893: out <= 16'h0532;    16'd43894: out <= 16'h0124;    16'd43895: out <= 16'h05A9;
    16'd43896: out <= 16'h002A;    16'd43897: out <= 16'h053C;    16'd43898: out <= 16'hFD0A;    16'd43899: out <= 16'h05C2;
    16'd43900: out <= 16'h0628;    16'd43901: out <= 16'hFB73;    16'd43902: out <= 16'h093F;    16'd43903: out <= 16'h09D3;
    16'd43904: out <= 16'h0461;    16'd43905: out <= 16'h03FA;    16'd43906: out <= 16'h0175;    16'd43907: out <= 16'h0141;
    16'd43908: out <= 16'h0A0F;    16'd43909: out <= 16'h029B;    16'd43910: out <= 16'h0294;    16'd43911: out <= 16'h079F;
    16'd43912: out <= 16'h0AEE;    16'd43913: out <= 16'h05F2;    16'd43914: out <= 16'h03B4;    16'd43915: out <= 16'hFD08;
    16'd43916: out <= 16'h05E7;    16'd43917: out <= 16'h0552;    16'd43918: out <= 16'h07A9;    16'd43919: out <= 16'h0192;
    16'd43920: out <= 16'h07F5;    16'd43921: out <= 16'h0898;    16'd43922: out <= 16'h03F1;    16'd43923: out <= 16'h0A54;
    16'd43924: out <= 16'h038E;    16'd43925: out <= 16'h0528;    16'd43926: out <= 16'h0602;    16'd43927: out <= 16'h019D;
    16'd43928: out <= 16'hFF27;    16'd43929: out <= 16'h0422;    16'd43930: out <= 16'h0458;    16'd43931: out <= 16'h0C32;
    16'd43932: out <= 16'h057A;    16'd43933: out <= 16'h04A4;    16'd43934: out <= 16'h054F;    16'd43935: out <= 16'h0746;
    16'd43936: out <= 16'h015C;    16'd43937: out <= 16'h0478;    16'd43938: out <= 16'h00A2;    16'd43939: out <= 16'h021F;
    16'd43940: out <= 16'h04BE;    16'd43941: out <= 16'h08CE;    16'd43942: out <= 16'h02F9;    16'd43943: out <= 16'h06BF;
    16'd43944: out <= 16'h001F;    16'd43945: out <= 16'h03CA;    16'd43946: out <= 16'h0032;    16'd43947: out <= 16'h019F;
    16'd43948: out <= 16'h0517;    16'd43949: out <= 16'h099A;    16'd43950: out <= 16'h0211;    16'd43951: out <= 16'h0583;
    16'd43952: out <= 16'h0394;    16'd43953: out <= 16'h057A;    16'd43954: out <= 16'hFF45;    16'd43955: out <= 16'h008A;
    16'd43956: out <= 16'h025B;    16'd43957: out <= 16'hFF08;    16'd43958: out <= 16'h002C;    16'd43959: out <= 16'h0187;
    16'd43960: out <= 16'h0627;    16'd43961: out <= 16'h03C2;    16'd43962: out <= 16'hFF6B;    16'd43963: out <= 16'h07C9;
    16'd43964: out <= 16'h0116;    16'd43965: out <= 16'h05B4;    16'd43966: out <= 16'h02A7;    16'd43967: out <= 16'h0644;
    16'd43968: out <= 16'h01E4;    16'd43969: out <= 16'h015D;    16'd43970: out <= 16'h0390;    16'd43971: out <= 16'h051A;
    16'd43972: out <= 16'h0756;    16'd43973: out <= 16'h0B5A;    16'd43974: out <= 16'h038B;    16'd43975: out <= 16'h09EA;
    16'd43976: out <= 16'h07A3;    16'd43977: out <= 16'h07AC;    16'd43978: out <= 16'h06B0;    16'd43979: out <= 16'h0800;
    16'd43980: out <= 16'hFFAA;    16'd43981: out <= 16'h042E;    16'd43982: out <= 16'h0A3E;    16'd43983: out <= 16'hFFCF;
    16'd43984: out <= 16'h01C6;    16'd43985: out <= 16'h06D2;    16'd43986: out <= 16'hFF3F;    16'd43987: out <= 16'hFE99;
    16'd43988: out <= 16'hFFD0;    16'd43989: out <= 16'h0579;    16'd43990: out <= 16'h06CB;    16'd43991: out <= 16'h05AF;
    16'd43992: out <= 16'hFAA7;    16'd43993: out <= 16'hFD01;    16'd43994: out <= 16'h0B75;    16'd43995: out <= 16'h002E;
    16'd43996: out <= 16'hFEEF;    16'd43997: out <= 16'hFD3C;    16'd43998: out <= 16'hFB01;    16'd43999: out <= 16'h0401;
    16'd44000: out <= 16'hF9B8;    16'd44001: out <= 16'hFBFA;    16'd44002: out <= 16'h041C;    16'd44003: out <= 16'h0331;
    16'd44004: out <= 16'h067D;    16'd44005: out <= 16'hFE3B;    16'd44006: out <= 16'h013C;    16'd44007: out <= 16'hFE12;
    16'd44008: out <= 16'h009C;    16'd44009: out <= 16'h03F3;    16'd44010: out <= 16'hFD36;    16'd44011: out <= 16'hFC74;
    16'd44012: out <= 16'h0123;    16'd44013: out <= 16'hFBB3;    16'd44014: out <= 16'hFE40;    16'd44015: out <= 16'h0847;
    16'd44016: out <= 16'h0191;    16'd44017: out <= 16'hF9DB;    16'd44018: out <= 16'h03CA;    16'd44019: out <= 16'hFDF5;
    16'd44020: out <= 16'h04CC;    16'd44021: out <= 16'hF8B8;    16'd44022: out <= 16'hFBE4;    16'd44023: out <= 16'hFDD9;
    16'd44024: out <= 16'h010A;    16'd44025: out <= 16'hFF4E;    16'd44026: out <= 16'h041D;    16'd44027: out <= 16'h0A73;
    16'd44028: out <= 16'hFDF5;    16'd44029: out <= 16'h0301;    16'd44030: out <= 16'hFB7E;    16'd44031: out <= 16'hFE5A;
    16'd44032: out <= 16'h0341;    16'd44033: out <= 16'h02D7;    16'd44034: out <= 16'hF86C;    16'd44035: out <= 16'hFFC7;
    16'd44036: out <= 16'h02E0;    16'd44037: out <= 16'hFF93;    16'd44038: out <= 16'h0511;    16'd44039: out <= 16'hFABC;
    16'd44040: out <= 16'hFD67;    16'd44041: out <= 16'h01D9;    16'd44042: out <= 16'h02D6;    16'd44043: out <= 16'h0041;
    16'd44044: out <= 16'hFC04;    16'd44045: out <= 16'h026F;    16'd44046: out <= 16'hF8E4;    16'd44047: out <= 16'h0330;
    16'd44048: out <= 16'h051F;    16'd44049: out <= 16'h03E8;    16'd44050: out <= 16'hFEA1;    16'd44051: out <= 16'hFCB6;
    16'd44052: out <= 16'h0050;    16'd44053: out <= 16'h04B5;    16'd44054: out <= 16'h0166;    16'd44055: out <= 16'h0013;
    16'd44056: out <= 16'h04F4;    16'd44057: out <= 16'h0267;    16'd44058: out <= 16'h02AD;    16'd44059: out <= 16'hFFD5;
    16'd44060: out <= 16'hFE20;    16'd44061: out <= 16'h03A3;    16'd44062: out <= 16'hFB38;    16'd44063: out <= 16'hFC12;
    16'd44064: out <= 16'h0353;    16'd44065: out <= 16'hFE26;    16'd44066: out <= 16'h0543;    16'd44067: out <= 16'h05D4;
    16'd44068: out <= 16'h09CC;    16'd44069: out <= 16'h018A;    16'd44070: out <= 16'h04A8;    16'd44071: out <= 16'h0454;
    16'd44072: out <= 16'h0838;    16'd44073: out <= 16'h00C1;    16'd44074: out <= 16'hFF26;    16'd44075: out <= 16'h021D;
    16'd44076: out <= 16'h0562;    16'd44077: out <= 16'h08D7;    16'd44078: out <= 16'hFF16;    16'd44079: out <= 16'h04AA;
    16'd44080: out <= 16'h054B;    16'd44081: out <= 16'h0692;    16'd44082: out <= 16'h0561;    16'd44083: out <= 16'h0037;
    16'd44084: out <= 16'h07C4;    16'd44085: out <= 16'hFF89;    16'd44086: out <= 16'h05AB;    16'd44087: out <= 16'h034A;
    16'd44088: out <= 16'h021F;    16'd44089: out <= 16'h0654;    16'd44090: out <= 16'h0464;    16'd44091: out <= 16'h07B3;
    16'd44092: out <= 16'h09A4;    16'd44093: out <= 16'h0C86;    16'd44094: out <= 16'h00BD;    16'd44095: out <= 16'h0748;
    16'd44096: out <= 16'h08E9;    16'd44097: out <= 16'h049B;    16'd44098: out <= 16'h07B0;    16'd44099: out <= 16'h020A;
    16'd44100: out <= 16'h01EA;    16'd44101: out <= 16'hFC4C;    16'd44102: out <= 16'h0155;    16'd44103: out <= 16'hFE63;
    16'd44104: out <= 16'h073E;    16'd44105: out <= 16'hFBE4;    16'd44106: out <= 16'h04E4;    16'd44107: out <= 16'h0D61;
    16'd44108: out <= 16'h034A;    16'd44109: out <= 16'h038F;    16'd44110: out <= 16'h07EA;    16'd44111: out <= 16'h033C;
    16'd44112: out <= 16'h044A;    16'd44113: out <= 16'h0495;    16'd44114: out <= 16'h0180;    16'd44115: out <= 16'hFFAF;
    16'd44116: out <= 16'h010A;    16'd44117: out <= 16'h0731;    16'd44118: out <= 16'h0A28;    16'd44119: out <= 16'h02AD;
    16'd44120: out <= 16'h0173;    16'd44121: out <= 16'h0018;    16'd44122: out <= 16'h03D9;    16'd44123: out <= 16'h0021;
    16'd44124: out <= 16'h068B;    16'd44125: out <= 16'h029C;    16'd44126: out <= 16'h0474;    16'd44127: out <= 16'h0054;
    16'd44128: out <= 16'h086B;    16'd44129: out <= 16'h02D9;    16'd44130: out <= 16'h0243;    16'd44131: out <= 16'h0716;
    16'd44132: out <= 16'h02ED;    16'd44133: out <= 16'h0101;    16'd44134: out <= 16'hFCE0;    16'd44135: out <= 16'hFEC8;
    16'd44136: out <= 16'h0385;    16'd44137: out <= 16'h0131;    16'd44138: out <= 16'h098C;    16'd44139: out <= 16'h01D6;
    16'd44140: out <= 16'h05CF;    16'd44141: out <= 16'h016F;    16'd44142: out <= 16'h0A09;    16'd44143: out <= 16'h092D;
    16'd44144: out <= 16'hFE26;    16'd44145: out <= 16'h029D;    16'd44146: out <= 16'hFE70;    16'd44147: out <= 16'h0635;
    16'd44148: out <= 16'h0607;    16'd44149: out <= 16'h0767;    16'd44150: out <= 16'h03E5;    16'd44151: out <= 16'h03EC;
    16'd44152: out <= 16'h0499;    16'd44153: out <= 16'h0068;    16'd44154: out <= 16'h023F;    16'd44155: out <= 16'h0391;
    16'd44156: out <= 16'h08EC;    16'd44157: out <= 16'h042E;    16'd44158: out <= 16'h023F;    16'd44159: out <= 16'h07AF;
    16'd44160: out <= 16'h0541;    16'd44161: out <= 16'h0644;    16'd44162: out <= 16'hFF80;    16'd44163: out <= 16'h055A;
    16'd44164: out <= 16'h0456;    16'd44165: out <= 16'h08B6;    16'd44166: out <= 16'h05D8;    16'd44167: out <= 16'h0586;
    16'd44168: out <= 16'hFF8E;    16'd44169: out <= 16'h00B0;    16'd44170: out <= 16'h035C;    16'd44171: out <= 16'h0447;
    16'd44172: out <= 16'h02E7;    16'd44173: out <= 16'h00E5;    16'd44174: out <= 16'h04EB;    16'd44175: out <= 16'h0555;
    16'd44176: out <= 16'hFF22;    16'd44177: out <= 16'h09E3;    16'd44178: out <= 16'h03BC;    16'd44179: out <= 16'h0392;
    16'd44180: out <= 16'h07ED;    16'd44181: out <= 16'h04A3;    16'd44182: out <= 16'h0328;    16'd44183: out <= 16'h03C6;
    16'd44184: out <= 16'h03B3;    16'd44185: out <= 16'h0043;    16'd44186: out <= 16'h0375;    16'd44187: out <= 16'h03E3;
    16'd44188: out <= 16'h096F;    16'd44189: out <= 16'h04B2;    16'd44190: out <= 16'hFE70;    16'd44191: out <= 16'h0840;
    16'd44192: out <= 16'hFCF1;    16'd44193: out <= 16'hFC1D;    16'd44194: out <= 16'h02AF;    16'd44195: out <= 16'h0ACF;
    16'd44196: out <= 16'hFC02;    16'd44197: out <= 16'h0A3B;    16'd44198: out <= 16'h01C1;    16'd44199: out <= 16'h0890;
    16'd44200: out <= 16'h0A4F;    16'd44201: out <= 16'h0276;    16'd44202: out <= 16'h006B;    16'd44203: out <= 16'h039D;
    16'd44204: out <= 16'h0CEA;    16'd44205: out <= 16'h0082;    16'd44206: out <= 16'hFF83;    16'd44207: out <= 16'h0738;
    16'd44208: out <= 16'h0ABA;    16'd44209: out <= 16'h07E5;    16'd44210: out <= 16'h0328;    16'd44211: out <= 16'h0191;
    16'd44212: out <= 16'h06E0;    16'd44213: out <= 16'hFF2D;    16'd44214: out <= 16'hF895;    16'd44215: out <= 16'h051D;
    16'd44216: out <= 16'h01A7;    16'd44217: out <= 16'h052B;    16'd44218: out <= 16'h0521;    16'd44219: out <= 16'h019A;
    16'd44220: out <= 16'h0379;    16'd44221: out <= 16'hFFE0;    16'd44222: out <= 16'h0222;    16'd44223: out <= 16'hFB3D;
    16'd44224: out <= 16'h04C5;    16'd44225: out <= 16'h004B;    16'd44226: out <= 16'h02ED;    16'd44227: out <= 16'h076B;
    16'd44228: out <= 16'h0516;    16'd44229: out <= 16'h0465;    16'd44230: out <= 16'hFFF8;    16'd44231: out <= 16'h0407;
    16'd44232: out <= 16'hFE16;    16'd44233: out <= 16'h00FF;    16'd44234: out <= 16'h0365;    16'd44235: out <= 16'h0039;
    16'd44236: out <= 16'h05BF;    16'd44237: out <= 16'h0BAD;    16'd44238: out <= 16'h0BB6;    16'd44239: out <= 16'h042B;
    16'd44240: out <= 16'h0492;    16'd44241: out <= 16'h0996;    16'd44242: out <= 16'h0A8B;    16'd44243: out <= 16'h0464;
    16'd44244: out <= 16'h054D;    16'd44245: out <= 16'h03B1;    16'd44246: out <= 16'h0340;    16'd44247: out <= 16'h00F9;
    16'd44248: out <= 16'h0245;    16'd44249: out <= 16'h0035;    16'd44250: out <= 16'hFF6F;    16'd44251: out <= 16'h0564;
    16'd44252: out <= 16'h074A;    16'd44253: out <= 16'hFF78;    16'd44254: out <= 16'h032B;    16'd44255: out <= 16'hFFF7;
    16'd44256: out <= 16'h039F;    16'd44257: out <= 16'h03E2;    16'd44258: out <= 16'h012A;    16'd44259: out <= 16'h0170;
    16'd44260: out <= 16'hFDB3;    16'd44261: out <= 16'hFD89;    16'd44262: out <= 16'h0370;    16'd44263: out <= 16'hFA1E;
    16'd44264: out <= 16'hFF6C;    16'd44265: out <= 16'h01E1;    16'd44266: out <= 16'h03FD;    16'd44267: out <= 16'hFFF6;
    16'd44268: out <= 16'h0128;    16'd44269: out <= 16'h04A4;    16'd44270: out <= 16'h09BC;    16'd44271: out <= 16'hFFB8;
    16'd44272: out <= 16'h04F3;    16'd44273: out <= 16'h006D;    16'd44274: out <= 16'h0176;    16'd44275: out <= 16'hFC65;
    16'd44276: out <= 16'hFB8C;    16'd44277: out <= 16'hFD3E;    16'd44278: out <= 16'h02BB;    16'd44279: out <= 16'hF972;
    16'd44280: out <= 16'h015C;    16'd44281: out <= 16'hFA71;    16'd44282: out <= 16'h01AB;    16'd44283: out <= 16'hF932;
    16'd44284: out <= 16'hF873;    16'd44285: out <= 16'h0535;    16'd44286: out <= 16'h0511;    16'd44287: out <= 16'h0293;
    16'd44288: out <= 16'h01B2;    16'd44289: out <= 16'hFF8E;    16'd44290: out <= 16'hFFA4;    16'd44291: out <= 16'h00A6;
    16'd44292: out <= 16'hF7DA;    16'd44293: out <= 16'h01C3;    16'd44294: out <= 16'hFD0B;    16'd44295: out <= 16'h0196;
    16'd44296: out <= 16'h0295;    16'd44297: out <= 16'hFFE7;    16'd44298: out <= 16'hFDD6;    16'd44299: out <= 16'h03BA;
    16'd44300: out <= 16'hFE8F;    16'd44301: out <= 16'h02AC;    16'd44302: out <= 16'hFF9B;    16'd44303: out <= 16'hFEA1;
    16'd44304: out <= 16'h048E;    16'd44305: out <= 16'hFDEF;    16'd44306: out <= 16'hFFFF;    16'd44307: out <= 16'hF68F;
    16'd44308: out <= 16'hFC3E;    16'd44309: out <= 16'h03C0;    16'd44310: out <= 16'h061F;    16'd44311: out <= 16'hFF0D;
    16'd44312: out <= 16'h00D6;    16'd44313: out <= 16'h067F;    16'd44314: out <= 16'h06E8;    16'd44315: out <= 16'h0384;
    16'd44316: out <= 16'hFFFF;    16'd44317: out <= 16'hFB4F;    16'd44318: out <= 16'hFE2A;    16'd44319: out <= 16'h04CA;
    16'd44320: out <= 16'h0172;    16'd44321: out <= 16'hF7D7;    16'd44322: out <= 16'h0161;    16'd44323: out <= 16'h08E6;
    16'd44324: out <= 16'h00D2;    16'd44325: out <= 16'h0064;    16'd44326: out <= 16'h097B;    16'd44327: out <= 16'h09DE;
    16'd44328: out <= 16'h0678;    16'd44329: out <= 16'h06B1;    16'd44330: out <= 16'hFFBD;    16'd44331: out <= 16'h0AF0;
    16'd44332: out <= 16'h031A;    16'd44333: out <= 16'h0C89;    16'd44334: out <= 16'h0276;    16'd44335: out <= 16'h0715;
    16'd44336: out <= 16'hFE74;    16'd44337: out <= 16'h0B63;    16'd44338: out <= 16'hFE40;    16'd44339: out <= 16'h0763;
    16'd44340: out <= 16'h072E;    16'd44341: out <= 16'h03FF;    16'd44342: out <= 16'h0250;    16'd44343: out <= 16'h00F9;
    16'd44344: out <= 16'h02D1;    16'd44345: out <= 16'h03D6;    16'd44346: out <= 16'h08E8;    16'd44347: out <= 16'h004D;
    16'd44348: out <= 16'h0698;    16'd44349: out <= 16'h0758;    16'd44350: out <= 16'h0704;    16'd44351: out <= 16'h0771;
    16'd44352: out <= 16'hFEE7;    16'd44353: out <= 16'h0471;    16'd44354: out <= 16'h02E9;    16'd44355: out <= 16'h0BC1;
    16'd44356: out <= 16'h03B1;    16'd44357: out <= 16'h00C3;    16'd44358: out <= 16'h0788;    16'd44359: out <= 16'h0631;
    16'd44360: out <= 16'h00CF;    16'd44361: out <= 16'hFF55;    16'd44362: out <= 16'h0208;    16'd44363: out <= 16'h07DB;
    16'd44364: out <= 16'hFD4A;    16'd44365: out <= 16'h0946;    16'd44366: out <= 16'h0834;    16'd44367: out <= 16'hFC57;
    16'd44368: out <= 16'h007C;    16'd44369: out <= 16'h05CC;    16'd44370: out <= 16'h06DF;    16'd44371: out <= 16'h0293;
    16'd44372: out <= 16'hFDCE;    16'd44373: out <= 16'h0633;    16'd44374: out <= 16'h0C38;    16'd44375: out <= 16'h011C;
    16'd44376: out <= 16'h0283;    16'd44377: out <= 16'h00F2;    16'd44378: out <= 16'h0576;    16'd44379: out <= 16'h02EF;
    16'd44380: out <= 16'h0013;    16'd44381: out <= 16'h0A65;    16'd44382: out <= 16'h062A;    16'd44383: out <= 16'h01F8;
    16'd44384: out <= 16'h04CD;    16'd44385: out <= 16'h053B;    16'd44386: out <= 16'h053D;    16'd44387: out <= 16'h0086;
    16'd44388: out <= 16'h0883;    16'd44389: out <= 16'h092F;    16'd44390: out <= 16'h0E00;    16'd44391: out <= 16'h0396;
    16'd44392: out <= 16'h004C;    16'd44393: out <= 16'hFD4E;    16'd44394: out <= 16'h0820;    16'd44395: out <= 16'h0192;
    16'd44396: out <= 16'hFD12;    16'd44397: out <= 16'h032A;    16'd44398: out <= 16'h03D6;    16'd44399: out <= 16'h0136;
    16'd44400: out <= 16'h0413;    16'd44401: out <= 16'h0921;    16'd44402: out <= 16'h0403;    16'd44403: out <= 16'h04C3;
    16'd44404: out <= 16'h0651;    16'd44405: out <= 16'h08B5;    16'd44406: out <= 16'h0261;    16'd44407: out <= 16'h05E2;
    16'd44408: out <= 16'h08EB;    16'd44409: out <= 16'h0401;    16'd44410: out <= 16'h0163;    16'd44411: out <= 16'h0574;
    16'd44412: out <= 16'h0578;    16'd44413: out <= 16'h0ACD;    16'd44414: out <= 16'h053A;    16'd44415: out <= 16'h05AE;
    16'd44416: out <= 16'h0A39;    16'd44417: out <= 16'hFED7;    16'd44418: out <= 16'h089D;    16'd44419: out <= 16'h03D2;
    16'd44420: out <= 16'h029E;    16'd44421: out <= 16'hFF1F;    16'd44422: out <= 16'h024D;    16'd44423: out <= 16'h08DA;
    16'd44424: out <= 16'h083F;    16'd44425: out <= 16'h04C4;    16'd44426: out <= 16'h0273;    16'd44427: out <= 16'h0054;
    16'd44428: out <= 16'hFDA0;    16'd44429: out <= 16'hFEC7;    16'd44430: out <= 16'hFED3;    16'd44431: out <= 16'h08F4;
    16'd44432: out <= 16'h084F;    16'd44433: out <= 16'h0389;    16'd44434: out <= 16'h02A8;    16'd44435: out <= 16'h09CC;
    16'd44436: out <= 16'h04A3;    16'd44437: out <= 16'h0702;    16'd44438: out <= 16'h02C2;    16'd44439: out <= 16'h0805;
    16'd44440: out <= 16'h026A;    16'd44441: out <= 16'h08C1;    16'd44442: out <= 16'h0596;    16'd44443: out <= 16'h0639;
    16'd44444: out <= 16'hFB3E;    16'd44445: out <= 16'h0210;    16'd44446: out <= 16'h0477;    16'd44447: out <= 16'hF9E5;
    16'd44448: out <= 16'hFF37;    16'd44449: out <= 16'h0598;    16'd44450: out <= 16'hFFD2;    16'd44451: out <= 16'h03F8;
    16'd44452: out <= 16'h08A7;    16'd44453: out <= 16'h0BD3;    16'd44454: out <= 16'h05E7;    16'd44455: out <= 16'h056C;
    16'd44456: out <= 16'h03DE;    16'd44457: out <= 16'h0401;    16'd44458: out <= 16'hFF9E;    16'd44459: out <= 16'hFFB1;
    16'd44460: out <= 16'h071A;    16'd44461: out <= 16'h016B;    16'd44462: out <= 16'h058A;    16'd44463: out <= 16'h02C4;
    16'd44464: out <= 16'h0084;    16'd44465: out <= 16'h07AA;    16'd44466: out <= 16'h01C7;    16'd44467: out <= 16'h0362;
    16'd44468: out <= 16'hFF43;    16'd44469: out <= 16'h00BE;    16'd44470: out <= 16'h02FF;    16'd44471: out <= 16'h0274;
    16'd44472: out <= 16'h00BD;    16'd44473: out <= 16'h07DE;    16'd44474: out <= 16'h04DE;    16'd44475: out <= 16'hFF06;
    16'd44476: out <= 16'h0C08;    16'd44477: out <= 16'h0129;    16'd44478: out <= 16'hFFCF;    16'd44479: out <= 16'h07CB;
    16'd44480: out <= 16'h000A;    16'd44481: out <= 16'hFF3D;    16'd44482: out <= 16'h01BC;    16'd44483: out <= 16'h0481;
    16'd44484: out <= 16'h0DD2;    16'd44485: out <= 16'h068A;    16'd44486: out <= 16'h0030;    16'd44487: out <= 16'h017A;
    16'd44488: out <= 16'h0234;    16'd44489: out <= 16'hFF4C;    16'd44490: out <= 16'h0823;    16'd44491: out <= 16'hFFB5;
    16'd44492: out <= 16'h02FA;    16'd44493: out <= 16'h005F;    16'd44494: out <= 16'h08E7;    16'd44495: out <= 16'h0329;
    16'd44496: out <= 16'h08C5;    16'd44497: out <= 16'h0830;    16'd44498: out <= 16'h0126;    16'd44499: out <= 16'h0510;
    16'd44500: out <= 16'h0613;    16'd44501: out <= 16'h06C3;    16'd44502: out <= 16'h0537;    16'd44503: out <= 16'hFCB7;
    16'd44504: out <= 16'hFF1C;    16'd44505: out <= 16'h00F5;    16'd44506: out <= 16'hFEED;    16'd44507: out <= 16'hFBCB;
    16'd44508: out <= 16'hFD37;    16'd44509: out <= 16'h0357;    16'd44510: out <= 16'h011C;    16'd44511: out <= 16'h0166;
    16'd44512: out <= 16'h02E7;    16'd44513: out <= 16'h0215;    16'd44514: out <= 16'h0244;    16'd44515: out <= 16'hFE21;
    16'd44516: out <= 16'hFBE1;    16'd44517: out <= 16'hFE34;    16'd44518: out <= 16'hFF48;    16'd44519: out <= 16'hFC46;
    16'd44520: out <= 16'hFC39;    16'd44521: out <= 16'hFCA3;    16'd44522: out <= 16'h0464;    16'd44523: out <= 16'h0172;
    16'd44524: out <= 16'h03AC;    16'd44525: out <= 16'h0410;    16'd44526: out <= 16'hFE99;    16'd44527: out <= 16'h0318;
    16'd44528: out <= 16'h0496;    16'd44529: out <= 16'hFAEC;    16'd44530: out <= 16'h05D4;    16'd44531: out <= 16'hFED3;
    16'd44532: out <= 16'hFDAC;    16'd44533: out <= 16'hFC3B;    16'd44534: out <= 16'h00F3;    16'd44535: out <= 16'h0104;
    16'd44536: out <= 16'hFF36;    16'd44537: out <= 16'h01F4;    16'd44538: out <= 16'hF3D5;    16'd44539: out <= 16'hFC83;
    16'd44540: out <= 16'h0483;    16'd44541: out <= 16'hFD7D;    16'd44542: out <= 16'hFFFA;    16'd44543: out <= 16'h02AE;
    16'd44544: out <= 16'hFBBC;    16'd44545: out <= 16'h00EE;    16'd44546: out <= 16'hFEBB;    16'd44547: out <= 16'h01EE;
    16'd44548: out <= 16'h0855;    16'd44549: out <= 16'hFCB4;    16'd44550: out <= 16'hFCD7;    16'd44551: out <= 16'hFDE0;
    16'd44552: out <= 16'hFD54;    16'd44553: out <= 16'hFA94;    16'd44554: out <= 16'h0207;    16'd44555: out <= 16'hF843;
    16'd44556: out <= 16'hF8B6;    16'd44557: out <= 16'hF8E1;    16'd44558: out <= 16'h04A9;    16'd44559: out <= 16'h043C;
    16'd44560: out <= 16'hFCC9;    16'd44561: out <= 16'hFF04;    16'd44562: out <= 16'h0207;    16'd44563: out <= 16'hFB0A;
    16'd44564: out <= 16'h098C;    16'd44565: out <= 16'hFE28;    16'd44566: out <= 16'hFB62;    16'd44567: out <= 16'h02CD;
    16'd44568: out <= 16'h01E6;    16'd44569: out <= 16'h02F4;    16'd44570: out <= 16'hFF83;    16'd44571: out <= 16'h06F8;
    16'd44572: out <= 16'hFECE;    16'd44573: out <= 16'hFDE2;    16'd44574: out <= 16'h0488;    16'd44575: out <= 16'h012E;
    16'd44576: out <= 16'hFE4D;    16'd44577: out <= 16'hFEB1;    16'd44578: out <= 16'h058F;    16'd44579: out <= 16'h048D;
    16'd44580: out <= 16'h014E;    16'd44581: out <= 16'h0E0E;    16'd44582: out <= 16'h073C;    16'd44583: out <= 16'h0037;
    16'd44584: out <= 16'h0540;    16'd44585: out <= 16'h032C;    16'd44586: out <= 16'h01A9;    16'd44587: out <= 16'hFE13;
    16'd44588: out <= 16'hFFFC;    16'd44589: out <= 16'hFEEA;    16'd44590: out <= 16'h050C;    16'd44591: out <= 16'h0406;
    16'd44592: out <= 16'h05C1;    16'd44593: out <= 16'h0C01;    16'd44594: out <= 16'h031F;    16'd44595: out <= 16'h03C9;
    16'd44596: out <= 16'h0254;    16'd44597: out <= 16'h02B1;    16'd44598: out <= 16'h00D6;    16'd44599: out <= 16'h04AA;
    16'd44600: out <= 16'h00CB;    16'd44601: out <= 16'h079B;    16'd44602: out <= 16'hFF66;    16'd44603: out <= 16'h078D;
    16'd44604: out <= 16'h0339;    16'd44605: out <= 16'h0496;    16'd44606: out <= 16'hFF42;    16'd44607: out <= 16'h08B5;
    16'd44608: out <= 16'h087E;    16'd44609: out <= 16'h0587;    16'd44610: out <= 16'h0593;    16'd44611: out <= 16'h0458;
    16'd44612: out <= 16'h010D;    16'd44613: out <= 16'h0ACE;    16'd44614: out <= 16'h0260;    16'd44615: out <= 16'h0450;
    16'd44616: out <= 16'hFEFB;    16'd44617: out <= 16'hFCE6;    16'd44618: out <= 16'h03B4;    16'd44619: out <= 16'h0867;
    16'd44620: out <= 16'h0130;    16'd44621: out <= 16'h044E;    16'd44622: out <= 16'h03A2;    16'd44623: out <= 16'h068D;
    16'd44624: out <= 16'h01DA;    16'd44625: out <= 16'hFBFE;    16'd44626: out <= 16'h060B;    16'd44627: out <= 16'h02B0;
    16'd44628: out <= 16'hFA2C;    16'd44629: out <= 16'hFC13;    16'd44630: out <= 16'h01F1;    16'd44631: out <= 16'hFCE0;
    16'd44632: out <= 16'h0367;    16'd44633: out <= 16'h05DD;    16'd44634: out <= 16'h0BA8;    16'd44635: out <= 16'h07CE;
    16'd44636: out <= 16'hFF74;    16'd44637: out <= 16'h00C7;    16'd44638: out <= 16'h0727;    16'd44639: out <= 16'h0439;
    16'd44640: out <= 16'h01A8;    16'd44641: out <= 16'h066F;    16'd44642: out <= 16'h0246;    16'd44643: out <= 16'hFE13;
    16'd44644: out <= 16'h0534;    16'd44645: out <= 16'h0028;    16'd44646: out <= 16'h0165;    16'd44647: out <= 16'h0997;
    16'd44648: out <= 16'h008F;    16'd44649: out <= 16'h0374;    16'd44650: out <= 16'h072E;    16'd44651: out <= 16'h0B53;
    16'd44652: out <= 16'h0085;    16'd44653: out <= 16'h034A;    16'd44654: out <= 16'hFFD1;    16'd44655: out <= 16'h04EC;
    16'd44656: out <= 16'h0145;    16'd44657: out <= 16'h0719;    16'd44658: out <= 16'h0B76;    16'd44659: out <= 16'h0183;
    16'd44660: out <= 16'h039D;    16'd44661: out <= 16'h0393;    16'd44662: out <= 16'h0810;    16'd44663: out <= 16'h0795;
    16'd44664: out <= 16'hF853;    16'd44665: out <= 16'hFF0F;    16'd44666: out <= 16'h0563;    16'd44667: out <= 16'h021C;
    16'd44668: out <= 16'hFFFF;    16'd44669: out <= 16'hFC46;    16'd44670: out <= 16'hFDF2;    16'd44671: out <= 16'h024D;
    16'd44672: out <= 16'h0676;    16'd44673: out <= 16'h0316;    16'd44674: out <= 16'h0574;    16'd44675: out <= 16'h0201;
    16'd44676: out <= 16'h04F3;    16'd44677: out <= 16'h064D;    16'd44678: out <= 16'h0183;    16'd44679: out <= 16'h01A4;
    16'd44680: out <= 16'h088C;    16'd44681: out <= 16'h05AF;    16'd44682: out <= 16'h0760;    16'd44683: out <= 16'h05C1;
    16'd44684: out <= 16'h003C;    16'd44685: out <= 16'h02AD;    16'd44686: out <= 16'h0A7A;    16'd44687: out <= 16'h0679;
    16'd44688: out <= 16'hFEA0;    16'd44689: out <= 16'hFFC2;    16'd44690: out <= 16'h09CD;    16'd44691: out <= 16'h0185;
    16'd44692: out <= 16'h012F;    16'd44693: out <= 16'hFA9A;    16'd44694: out <= 16'h091A;    16'd44695: out <= 16'h0735;
    16'd44696: out <= 16'hFADF;    16'd44697: out <= 16'h0621;    16'd44698: out <= 16'h07EF;    16'd44699: out <= 16'hFDAC;
    16'd44700: out <= 16'h0A5C;    16'd44701: out <= 16'h02FE;    16'd44702: out <= 16'h02FC;    16'd44703: out <= 16'hFC68;
    16'd44704: out <= 16'h0576;    16'd44705: out <= 16'h0875;    16'd44706: out <= 16'h04D1;    16'd44707: out <= 16'h01ED;
    16'd44708: out <= 16'hF833;    16'd44709: out <= 16'h094F;    16'd44710: out <= 16'h05B8;    16'd44711: out <= 16'h082A;
    16'd44712: out <= 16'hFD32;    16'd44713: out <= 16'hFDA5;    16'd44714: out <= 16'h0544;    16'd44715: out <= 16'h0C8E;
    16'd44716: out <= 16'h09C3;    16'd44717: out <= 16'h07EB;    16'd44718: out <= 16'h00E6;    16'd44719: out <= 16'h08C4;
    16'd44720: out <= 16'h07A4;    16'd44721: out <= 16'h0359;    16'd44722: out <= 16'h070D;    16'd44723: out <= 16'h0417;
    16'd44724: out <= 16'h0589;    16'd44725: out <= 16'h042B;    16'd44726: out <= 16'h0404;    16'd44727: out <= 16'h0716;
    16'd44728: out <= 16'h06EF;    16'd44729: out <= 16'h010C;    16'd44730: out <= 16'h0361;    16'd44731: out <= 16'h00A4;
    16'd44732: out <= 16'h07C4;    16'd44733: out <= 16'h0167;    16'd44734: out <= 16'h0D31;    16'd44735: out <= 16'h0357;
    16'd44736: out <= 16'h029C;    16'd44737: out <= 16'h0101;    16'd44738: out <= 16'h05D9;    16'd44739: out <= 16'h04DC;
    16'd44740: out <= 16'h03A0;    16'd44741: out <= 16'hFFDF;    16'd44742: out <= 16'h04A1;    16'd44743: out <= 16'h04B9;
    16'd44744: out <= 16'h0136;    16'd44745: out <= 16'h0624;    16'd44746: out <= 16'hFDB1;    16'd44747: out <= 16'h026F;
    16'd44748: out <= 16'h0119;    16'd44749: out <= 16'hFD57;    16'd44750: out <= 16'hFDAB;    16'd44751: out <= 16'hF9E4;
    16'd44752: out <= 16'h0647;    16'd44753: out <= 16'hFEAF;    16'd44754: out <= 16'hFA53;    16'd44755: out <= 16'h045C;
    16'd44756: out <= 16'hFB05;    16'd44757: out <= 16'hFB2E;    16'd44758: out <= 16'h0029;    16'd44759: out <= 16'hFCB8;
    16'd44760: out <= 16'h044C;    16'd44761: out <= 16'h025E;    16'd44762: out <= 16'h0024;    16'd44763: out <= 16'hFA9C;
    16'd44764: out <= 16'h0137;    16'd44765: out <= 16'hFCFC;    16'd44766: out <= 16'hFA78;    16'd44767: out <= 16'h05D3;
    16'd44768: out <= 16'h037A;    16'd44769: out <= 16'hFFDD;    16'd44770: out <= 16'h040C;    16'd44771: out <= 16'hFFDA;
    16'd44772: out <= 16'h036E;    16'd44773: out <= 16'hFEB4;    16'd44774: out <= 16'hFA64;    16'd44775: out <= 16'h0256;
    16'd44776: out <= 16'hFE79;    16'd44777: out <= 16'hFE28;    16'd44778: out <= 16'h009F;    16'd44779: out <= 16'h04D3;
    16'd44780: out <= 16'h01A7;    16'd44781: out <= 16'h017E;    16'd44782: out <= 16'hFE6B;    16'd44783: out <= 16'h0532;
    16'd44784: out <= 16'h01F6;    16'd44785: out <= 16'h05BD;    16'd44786: out <= 16'hFC98;    16'd44787: out <= 16'h040A;
    16'd44788: out <= 16'h027E;    16'd44789: out <= 16'h0010;    16'd44790: out <= 16'h04B3;    16'd44791: out <= 16'h0651;
    16'd44792: out <= 16'h02A1;    16'd44793: out <= 16'hFC5F;    16'd44794: out <= 16'hFF90;    16'd44795: out <= 16'hFB70;
    16'd44796: out <= 16'hFC02;    16'd44797: out <= 16'hFB72;    16'd44798: out <= 16'h0238;    16'd44799: out <= 16'hFE5B;
    16'd44800: out <= 16'h00E0;    16'd44801: out <= 16'h02A6;    16'd44802: out <= 16'h01DC;    16'd44803: out <= 16'hF95E;
    16'd44804: out <= 16'h04E4;    16'd44805: out <= 16'h020E;    16'd44806: out <= 16'h0344;    16'd44807: out <= 16'hFB13;
    16'd44808: out <= 16'hFC60;    16'd44809: out <= 16'h06CC;    16'd44810: out <= 16'hFE46;    16'd44811: out <= 16'hFBEF;
    16'd44812: out <= 16'h005A;    16'd44813: out <= 16'hFAE9;    16'd44814: out <= 16'h002F;    16'd44815: out <= 16'hFD95;
    16'd44816: out <= 16'hFC7A;    16'd44817: out <= 16'hFC46;    16'd44818: out <= 16'h016F;    16'd44819: out <= 16'h0301;
    16'd44820: out <= 16'hFFE3;    16'd44821: out <= 16'h02D7;    16'd44822: out <= 16'h0184;    16'd44823: out <= 16'hFE89;
    16'd44824: out <= 16'hFE2B;    16'd44825: out <= 16'hFB06;    16'd44826: out <= 16'hFC3D;    16'd44827: out <= 16'h0202;
    16'd44828: out <= 16'h0643;    16'd44829: out <= 16'hFB0B;    16'd44830: out <= 16'h02C8;    16'd44831: out <= 16'hFC42;
    16'd44832: out <= 16'h0001;    16'd44833: out <= 16'h01C3;    16'd44834: out <= 16'h0189;    16'd44835: out <= 16'h02C1;
    16'd44836: out <= 16'h0E2A;    16'd44837: out <= 16'h06CB;    16'd44838: out <= 16'h0167;    16'd44839: out <= 16'hFE96;
    16'd44840: out <= 16'h02C9;    16'd44841: out <= 16'hFDC1;    16'd44842: out <= 16'h072A;    16'd44843: out <= 16'h04CD;
    16'd44844: out <= 16'h0595;    16'd44845: out <= 16'h03C0;    16'd44846: out <= 16'h047D;    16'd44847: out <= 16'h0396;
    16'd44848: out <= 16'h05B5;    16'd44849: out <= 16'h02A5;    16'd44850: out <= 16'h02BD;    16'd44851: out <= 16'h01E0;
    16'd44852: out <= 16'hFFC4;    16'd44853: out <= 16'h0787;    16'd44854: out <= 16'hFE2F;    16'd44855: out <= 16'h04C7;
    16'd44856: out <= 16'h0787;    16'd44857: out <= 16'h0067;    16'd44858: out <= 16'h05A4;    16'd44859: out <= 16'hFAC9;
    16'd44860: out <= 16'h02BD;    16'd44861: out <= 16'h03A9;    16'd44862: out <= 16'h03A8;    16'd44863: out <= 16'h0254;
    16'd44864: out <= 16'h055A;    16'd44865: out <= 16'h04B2;    16'd44866: out <= 16'h057D;    16'd44867: out <= 16'h0954;
    16'd44868: out <= 16'hFF48;    16'd44869: out <= 16'h057E;    16'd44870: out <= 16'h0481;    16'd44871: out <= 16'h02F0;
    16'd44872: out <= 16'h0945;    16'd44873: out <= 16'hFDC9;    16'd44874: out <= 16'h0673;    16'd44875: out <= 16'h038D;
    16'd44876: out <= 16'h067A;    16'd44877: out <= 16'hFDF1;    16'd44878: out <= 16'h04B7;    16'd44879: out <= 16'h02FE;
    16'd44880: out <= 16'h04ED;    16'd44881: out <= 16'h04B6;    16'd44882: out <= 16'h05C8;    16'd44883: out <= 16'h03A6;
    16'd44884: out <= 16'h073C;    16'd44885: out <= 16'h00B9;    16'd44886: out <= 16'h080F;    16'd44887: out <= 16'h02E4;
    16'd44888: out <= 16'h001E;    16'd44889: out <= 16'hFFF6;    16'd44890: out <= 16'h008F;    16'd44891: out <= 16'h04D8;
    16'd44892: out <= 16'h0885;    16'd44893: out <= 16'h026B;    16'd44894: out <= 16'h0693;    16'd44895: out <= 16'hF780;
    16'd44896: out <= 16'h0882;    16'd44897: out <= 16'h0A4C;    16'd44898: out <= 16'h09B3;    16'd44899: out <= 16'hFFD4;
    16'd44900: out <= 16'h00F1;    16'd44901: out <= 16'h0356;    16'd44902: out <= 16'h01D2;    16'd44903: out <= 16'h0878;
    16'd44904: out <= 16'h0049;    16'd44905: out <= 16'h06C0;    16'd44906: out <= 16'h082D;    16'd44907: out <= 16'h03A3;
    16'd44908: out <= 16'h090F;    16'd44909: out <= 16'h0739;    16'd44910: out <= 16'h0204;    16'd44911: out <= 16'h058B;
    16'd44912: out <= 16'h01A4;    16'd44913: out <= 16'h02A9;    16'd44914: out <= 16'h0327;    16'd44915: out <= 16'h0528;
    16'd44916: out <= 16'h0932;    16'd44917: out <= 16'h0A96;    16'd44918: out <= 16'h0789;    16'd44919: out <= 16'h0742;
    16'd44920: out <= 16'h00A2;    16'd44921: out <= 16'h0744;    16'd44922: out <= 16'h03A5;    16'd44923: out <= 16'h073E;
    16'd44924: out <= 16'hFEB9;    16'd44925: out <= 16'h049D;    16'd44926: out <= 16'h059D;    16'd44927: out <= 16'h0748;
    16'd44928: out <= 16'h07F3;    16'd44929: out <= 16'h0455;    16'd44930: out <= 16'h054C;    16'd44931: out <= 16'h04E0;
    16'd44932: out <= 16'h0340;    16'd44933: out <= 16'h00A8;    16'd44934: out <= 16'h0933;    16'd44935: out <= 16'h048F;
    16'd44936: out <= 16'h031D;    16'd44937: out <= 16'h008E;    16'd44938: out <= 16'h0271;    16'd44939: out <= 16'h02AD;
    16'd44940: out <= 16'h05AD;    16'd44941: out <= 16'h03CF;    16'd44942: out <= 16'h03C4;    16'd44943: out <= 16'hFFAF;
    16'd44944: out <= 16'h0281;    16'd44945: out <= 16'h0A1F;    16'd44946: out <= 16'h0276;    16'd44947: out <= 16'h07D8;
    16'd44948: out <= 16'h005B;    16'd44949: out <= 16'h0532;    16'd44950: out <= 16'h015E;    16'd44951: out <= 16'hFEBB;
    16'd44952: out <= 16'h0710;    16'd44953: out <= 16'h055E;    16'd44954: out <= 16'hFCB1;    16'd44955: out <= 16'h04E9;
    16'd44956: out <= 16'h031D;    16'd44957: out <= 16'h0646;    16'd44958: out <= 16'hFC25;    16'd44959: out <= 16'h0342;
    16'd44960: out <= 16'hF8EA;    16'd44961: out <= 16'h03F5;    16'd44962: out <= 16'h003A;    16'd44963: out <= 16'h0328;
    16'd44964: out <= 16'hFC0A;    16'd44965: out <= 16'h06E7;    16'd44966: out <= 16'h024A;    16'd44967: out <= 16'h059C;
    16'd44968: out <= 16'h0BC8;    16'd44969: out <= 16'h01E7;    16'd44970: out <= 16'h00AB;    16'd44971: out <= 16'hFF46;
    16'd44972: out <= 16'h00C5;    16'd44973: out <= 16'h022E;    16'd44974: out <= 16'h00D0;    16'd44975: out <= 16'h05A2;
    16'd44976: out <= 16'h038C;    16'd44977: out <= 16'h053E;    16'd44978: out <= 16'hFF3B;    16'd44979: out <= 16'h058E;
    16'd44980: out <= 16'h0119;    16'd44981: out <= 16'hFE6B;    16'd44982: out <= 16'h016F;    16'd44983: out <= 16'hFD7C;
    16'd44984: out <= 16'hFEF1;    16'd44985: out <= 16'h0923;    16'd44986: out <= 16'h07E2;    16'd44987: out <= 16'h02E1;
    16'd44988: out <= 16'h0041;    16'd44989: out <= 16'h07ED;    16'd44990: out <= 16'h02CF;    16'd44991: out <= 16'hFF4D;
    16'd44992: out <= 16'h0241;    16'd44993: out <= 16'h06A8;    16'd44994: out <= 16'h0697;    16'd44995: out <= 16'h091C;
    16'd44996: out <= 16'h0742;    16'd44997: out <= 16'hFC95;    16'd44998: out <= 16'h020B;    16'd44999: out <= 16'h091B;
    16'd45000: out <= 16'h06EB;    16'd45001: out <= 16'h022A;    16'd45002: out <= 16'h034B;    16'd45003: out <= 16'h0043;
    16'd45004: out <= 16'h0103;    16'd45005: out <= 16'hFF02;    16'd45006: out <= 16'h05F5;    16'd45007: out <= 16'hFBC7;
    16'd45008: out <= 16'hFEB4;    16'd45009: out <= 16'hFC3D;    16'd45010: out <= 16'h01BB;    16'd45011: out <= 16'h0311;
    16'd45012: out <= 16'hF6EB;    16'd45013: out <= 16'h013D;    16'd45014: out <= 16'h0381;    16'd45015: out <= 16'hFEA5;
    16'd45016: out <= 16'hFEC1;    16'd45017: out <= 16'h087D;    16'd45018: out <= 16'hF74A;    16'd45019: out <= 16'hFEEF;
    16'd45020: out <= 16'hF9CD;    16'd45021: out <= 16'h002D;    16'd45022: out <= 16'h031E;    16'd45023: out <= 16'hFE7A;
    16'd45024: out <= 16'hF956;    16'd45025: out <= 16'hFE3E;    16'd45026: out <= 16'hFF6C;    16'd45027: out <= 16'hFBE6;
    16'd45028: out <= 16'h0358;    16'd45029: out <= 16'h004F;    16'd45030: out <= 16'h031C;    16'd45031: out <= 16'hFB8C;
    16'd45032: out <= 16'hFB7C;    16'd45033: out <= 16'hFE65;    16'd45034: out <= 16'h0050;    16'd45035: out <= 16'hFEFC;
    16'd45036: out <= 16'hFF9E;    16'd45037: out <= 16'hFEDA;    16'd45038: out <= 16'hFFE7;    16'd45039: out <= 16'h0441;
    16'd45040: out <= 16'h068E;    16'd45041: out <= 16'h021C;    16'd45042: out <= 16'hFF03;    16'd45043: out <= 16'hFCE8;
    16'd45044: out <= 16'hFC41;    16'd45045: out <= 16'hFF1E;    16'd45046: out <= 16'hFF5E;    16'd45047: out <= 16'h0265;
    16'd45048: out <= 16'hFEDA;    16'd45049: out <= 16'hFAE2;    16'd45050: out <= 16'hFB09;    16'd45051: out <= 16'hFC4B;
    16'd45052: out <= 16'hFE03;    16'd45053: out <= 16'hFFFB;    16'd45054: out <= 16'hFDC4;    16'd45055: out <= 16'h03AA;
    16'd45056: out <= 16'h010B;    16'd45057: out <= 16'h012E;    16'd45058: out <= 16'hFC7A;    16'd45059: out <= 16'h03F1;
    16'd45060: out <= 16'hFFBB;    16'd45061: out <= 16'h013E;    16'd45062: out <= 16'h01ED;    16'd45063: out <= 16'h0090;
    16'd45064: out <= 16'hFBB9;    16'd45065: out <= 16'h01C6;    16'd45066: out <= 16'h0436;    16'd45067: out <= 16'hFEF9;
    16'd45068: out <= 16'hFE3F;    16'd45069: out <= 16'hFEF3;    16'd45070: out <= 16'h00B8;    16'd45071: out <= 16'h028B;
    16'd45072: out <= 16'hFE9C;    16'd45073: out <= 16'hF846;    16'd45074: out <= 16'h002D;    16'd45075: out <= 16'hFE1B;
    16'd45076: out <= 16'hFFB8;    16'd45077: out <= 16'hFEC8;    16'd45078: out <= 16'h05FF;    16'd45079: out <= 16'hFEF9;
    16'd45080: out <= 16'hFF87;    16'd45081: out <= 16'h0838;    16'd45082: out <= 16'hFCF9;    16'd45083: out <= 16'hF94A;
    16'd45084: out <= 16'h0170;    16'd45085: out <= 16'hFAB3;    16'd45086: out <= 16'h0846;    16'd45087: out <= 16'h0201;
    16'd45088: out <= 16'hFE01;    16'd45089: out <= 16'h0815;    16'd45090: out <= 16'h000A;    16'd45091: out <= 16'h09CC;
    16'd45092: out <= 16'hFAC3;    16'd45093: out <= 16'h0302;    16'd45094: out <= 16'h095C;    16'd45095: out <= 16'h0446;
    16'd45096: out <= 16'h005A;    16'd45097: out <= 16'h0163;    16'd45098: out <= 16'h050D;    16'd45099: out <= 16'h03C4;
    16'd45100: out <= 16'h0BE4;    16'd45101: out <= 16'h0373;    16'd45102: out <= 16'h00C7;    16'd45103: out <= 16'h0482;
    16'd45104: out <= 16'h02C7;    16'd45105: out <= 16'h023C;    16'd45106: out <= 16'h0A20;    16'd45107: out <= 16'h024A;
    16'd45108: out <= 16'h045D;    16'd45109: out <= 16'hFA68;    16'd45110: out <= 16'h02C4;    16'd45111: out <= 16'h061F;
    16'd45112: out <= 16'hFD67;    16'd45113: out <= 16'h0A44;    16'd45114: out <= 16'h0ED2;    16'd45115: out <= 16'hFC90;
    16'd45116: out <= 16'h0581;    16'd45117: out <= 16'h0A01;    16'd45118: out <= 16'h0305;    16'd45119: out <= 16'h09B7;
    16'd45120: out <= 16'h0710;    16'd45121: out <= 16'h007C;    16'd45122: out <= 16'h01EF;    16'd45123: out <= 16'h05A3;
    16'd45124: out <= 16'h084D;    16'd45125: out <= 16'h0341;    16'd45126: out <= 16'h041E;    16'd45127: out <= 16'h07B4;
    16'd45128: out <= 16'h04F3;    16'd45129: out <= 16'hFFBD;    16'd45130: out <= 16'h047A;    16'd45131: out <= 16'h0738;
    16'd45132: out <= 16'h021B;    16'd45133: out <= 16'h06AC;    16'd45134: out <= 16'h06E9;    16'd45135: out <= 16'h0BB5;
    16'd45136: out <= 16'h08D3;    16'd45137: out <= 16'h02AA;    16'd45138: out <= 16'h05AE;    16'd45139: out <= 16'h045D;
    16'd45140: out <= 16'h01C8;    16'd45141: out <= 16'h04F5;    16'd45142: out <= 16'h0E9D;    16'd45143: out <= 16'h03E1;
    16'd45144: out <= 16'h0432;    16'd45145: out <= 16'h04A2;    16'd45146: out <= 16'h00BD;    16'd45147: out <= 16'h00A9;
    16'd45148: out <= 16'h0498;    16'd45149: out <= 16'h0AC3;    16'd45150: out <= 16'h062C;    16'd45151: out <= 16'h0337;
    16'd45152: out <= 16'hFD30;    16'd45153: out <= 16'h00A8;    16'd45154: out <= 16'h093B;    16'd45155: out <= 16'h0890;
    16'd45156: out <= 16'h08DA;    16'd45157: out <= 16'h05A9;    16'd45158: out <= 16'hFE3E;    16'd45159: out <= 16'h0543;
    16'd45160: out <= 16'h059C;    16'd45161: out <= 16'h061A;    16'd45162: out <= 16'hFFB3;    16'd45163: out <= 16'h0B0D;
    16'd45164: out <= 16'h0C0F;    16'd45165: out <= 16'hFBB3;    16'd45166: out <= 16'hFFCD;    16'd45167: out <= 16'hFB2E;
    16'd45168: out <= 16'h028C;    16'd45169: out <= 16'h0247;    16'd45170: out <= 16'hFF97;    16'd45171: out <= 16'hF825;
    16'd45172: out <= 16'h00F4;    16'd45173: out <= 16'h0529;    16'd45174: out <= 16'h029D;    16'd45175: out <= 16'hFAF1;
    16'd45176: out <= 16'h0632;    16'd45177: out <= 16'h072C;    16'd45178: out <= 16'h01A2;    16'd45179: out <= 16'h026A;
    16'd45180: out <= 16'h0086;    16'd45181: out <= 16'h02F0;    16'd45182: out <= 16'h0239;    16'd45183: out <= 16'h0640;
    16'd45184: out <= 16'hFE5A;    16'd45185: out <= 16'h01DC;    16'd45186: out <= 16'h0476;    16'd45187: out <= 16'hFB6B;
    16'd45188: out <= 16'h0634;    16'd45189: out <= 16'h03BC;    16'd45190: out <= 16'hFF66;    16'd45191: out <= 16'h0382;
    16'd45192: out <= 16'h05C3;    16'd45193: out <= 16'h0753;    16'd45194: out <= 16'h0328;    16'd45195: out <= 16'h0127;
    16'd45196: out <= 16'h0321;    16'd45197: out <= 16'h03A0;    16'd45198: out <= 16'h012F;    16'd45199: out <= 16'h03DF;
    16'd45200: out <= 16'h0253;    16'd45201: out <= 16'hFB87;    16'd45202: out <= 16'h048D;    16'd45203: out <= 16'h052D;
    16'd45204: out <= 16'h0495;    16'd45205: out <= 16'h0360;    16'd45206: out <= 16'h0337;    16'd45207: out <= 16'h091C;
    16'd45208: out <= 16'h04C5;    16'd45209: out <= 16'h01E5;    16'd45210: out <= 16'hFF8D;    16'd45211: out <= 16'h07CA;
    16'd45212: out <= 16'h0478;    16'd45213: out <= 16'h0C8E;    16'd45214: out <= 16'h07DA;    16'd45215: out <= 16'h055C;
    16'd45216: out <= 16'h033B;    16'd45217: out <= 16'h05E8;    16'd45218: out <= 16'h00C2;    16'd45219: out <= 16'h059E;
    16'd45220: out <= 16'h007D;    16'd45221: out <= 16'h043F;    16'd45222: out <= 16'h0551;    16'd45223: out <= 16'h04A5;
    16'd45224: out <= 16'h095B;    16'd45225: out <= 16'h050A;    16'd45226: out <= 16'h0287;    16'd45227: out <= 16'h0229;
    16'd45228: out <= 16'h033A;    16'd45229: out <= 16'h002A;    16'd45230: out <= 16'hFD6C;    16'd45231: out <= 16'h045C;
    16'd45232: out <= 16'h02C7;    16'd45233: out <= 16'h00C8;    16'd45234: out <= 16'h091C;    16'd45235: out <= 16'h079B;
    16'd45236: out <= 16'h00DF;    16'd45237: out <= 16'h03EA;    16'd45238: out <= 16'h0216;    16'd45239: out <= 16'h021B;
    16'd45240: out <= 16'h06EF;    16'd45241: out <= 16'h00F6;    16'd45242: out <= 16'h039D;    16'd45243: out <= 16'h0305;
    16'd45244: out <= 16'hFE6B;    16'd45245: out <= 16'h0754;    16'd45246: out <= 16'h04F6;    16'd45247: out <= 16'h0230;
    16'd45248: out <= 16'h016E;    16'd45249: out <= 16'h007A;    16'd45250: out <= 16'h01B0;    16'd45251: out <= 16'h0381;
    16'd45252: out <= 16'h0BF6;    16'd45253: out <= 16'h00EE;    16'd45254: out <= 16'h08C4;    16'd45255: out <= 16'h064B;
    16'd45256: out <= 16'h04E0;    16'd45257: out <= 16'h05F7;    16'd45258: out <= 16'h09D0;    16'd45259: out <= 16'h0045;
    16'd45260: out <= 16'h07D7;    16'd45261: out <= 16'h049B;    16'd45262: out <= 16'hFD6F;    16'd45263: out <= 16'hFC2D;
    16'd45264: out <= 16'h02B6;    16'd45265: out <= 16'hFD36;    16'd45266: out <= 16'h0518;    16'd45267: out <= 16'h025C;
    16'd45268: out <= 16'hFA40;    16'd45269: out <= 16'hFCBA;    16'd45270: out <= 16'h013D;    16'd45271: out <= 16'hFEEF;
    16'd45272: out <= 16'h00C2;    16'd45273: out <= 16'h047B;    16'd45274: out <= 16'hFE90;    16'd45275: out <= 16'h018D;
    16'd45276: out <= 16'hFA03;    16'd45277: out <= 16'hFF8D;    16'd45278: out <= 16'hFD96;    16'd45279: out <= 16'h0287;
    16'd45280: out <= 16'h036B;    16'd45281: out <= 16'h0177;    16'd45282: out <= 16'hFDDF;    16'd45283: out <= 16'h01E3;
    16'd45284: out <= 16'h020A;    16'd45285: out <= 16'h0739;    16'd45286: out <= 16'hFD02;    16'd45287: out <= 16'hFB67;
    16'd45288: out <= 16'h00BB;    16'd45289: out <= 16'h028A;    16'd45290: out <= 16'h006B;    16'd45291: out <= 16'hF5BE;
    16'd45292: out <= 16'h04AC;    16'd45293: out <= 16'hFD81;    16'd45294: out <= 16'hF971;    16'd45295: out <= 16'h01B0;
    16'd45296: out <= 16'hFA57;    16'd45297: out <= 16'h0431;    16'd45298: out <= 16'h0313;    16'd45299: out <= 16'h0260;
    16'd45300: out <= 16'hFDB6;    16'd45301: out <= 16'hFBD6;    16'd45302: out <= 16'hFCA3;    16'd45303: out <= 16'hFD67;
    16'd45304: out <= 16'hFE1D;    16'd45305: out <= 16'h00C0;    16'd45306: out <= 16'h019B;    16'd45307: out <= 16'h009A;
    16'd45308: out <= 16'h0387;    16'd45309: out <= 16'hFB68;    16'd45310: out <= 16'h020B;    16'd45311: out <= 16'h01BE;
    16'd45312: out <= 16'h095F;    16'd45313: out <= 16'h061B;    16'd45314: out <= 16'h004A;    16'd45315: out <= 16'hF7B5;
    16'd45316: out <= 16'h00FD;    16'd45317: out <= 16'hFFF1;    16'd45318: out <= 16'h057F;    16'd45319: out <= 16'hFF15;
    16'd45320: out <= 16'h0056;    16'd45321: out <= 16'hFC44;    16'd45322: out <= 16'h010F;    16'd45323: out <= 16'hFABB;
    16'd45324: out <= 16'hF805;    16'd45325: out <= 16'hFD90;    16'd45326: out <= 16'h02FD;    16'd45327: out <= 16'h01B4;
    16'd45328: out <= 16'h0461;    16'd45329: out <= 16'h02BC;    16'd45330: out <= 16'hFE56;    16'd45331: out <= 16'hFC47;
    16'd45332: out <= 16'h00E5;    16'd45333: out <= 16'h00F1;    16'd45334: out <= 16'h04B7;    16'd45335: out <= 16'hFFDF;
    16'd45336: out <= 16'h02E8;    16'd45337: out <= 16'hFE0B;    16'd45338: out <= 16'h016A;    16'd45339: out <= 16'hFB21;
    16'd45340: out <= 16'h01E5;    16'd45341: out <= 16'h01C9;    16'd45342: out <= 16'h00C2;    16'd45343: out <= 16'hF85A;
    16'd45344: out <= 16'hFF77;    16'd45345: out <= 16'hFF12;    16'd45346: out <= 16'hFD3D;    16'd45347: out <= 16'hFE15;
    16'd45348: out <= 16'h0881;    16'd45349: out <= 16'h0B51;    16'd45350: out <= 16'hFF11;    16'd45351: out <= 16'h00E0;
    16'd45352: out <= 16'hFC4A;    16'd45353: out <= 16'h0080;    16'd45354: out <= 16'h04D1;    16'd45355: out <= 16'h018B;
    16'd45356: out <= 16'h0276;    16'd45357: out <= 16'h0586;    16'd45358: out <= 16'h0497;    16'd45359: out <= 16'h06C8;
    16'd45360: out <= 16'h0209;    16'd45361: out <= 16'hFE41;    16'd45362: out <= 16'h0287;    16'd45363: out <= 16'h01FB;
    16'd45364: out <= 16'h0357;    16'd45365: out <= 16'h04F6;    16'd45366: out <= 16'h053C;    16'd45367: out <= 16'h01EC;
    16'd45368: out <= 16'h0776;    16'd45369: out <= 16'h062C;    16'd45370: out <= 16'h01C5;    16'd45371: out <= 16'h0132;
    16'd45372: out <= 16'h0296;    16'd45373: out <= 16'h0726;    16'd45374: out <= 16'h0348;    16'd45375: out <= 16'h0786;
    16'd45376: out <= 16'h059A;    16'd45377: out <= 16'h0663;    16'd45378: out <= 16'h05E7;    16'd45379: out <= 16'h085B;
    16'd45380: out <= 16'h08C5;    16'd45381: out <= 16'h0692;    16'd45382: out <= 16'h0770;    16'd45383: out <= 16'h0829;
    16'd45384: out <= 16'h0006;    16'd45385: out <= 16'h048C;    16'd45386: out <= 16'h03EB;    16'd45387: out <= 16'h0589;
    16'd45388: out <= 16'h0847;    16'd45389: out <= 16'h0172;    16'd45390: out <= 16'h05D4;    16'd45391: out <= 16'h032B;
    16'd45392: out <= 16'h02BE;    16'd45393: out <= 16'h004C;    16'd45394: out <= 16'h05EF;    16'd45395: out <= 16'h00E8;
    16'd45396: out <= 16'hFF0B;    16'd45397: out <= 16'hFF7B;    16'd45398: out <= 16'h00EB;    16'd45399: out <= 16'h056A;
    16'd45400: out <= 16'h07A3;    16'd45401: out <= 16'hFBC8;    16'd45402: out <= 16'h0A69;    16'd45403: out <= 16'h05AA;
    16'd45404: out <= 16'h046B;    16'd45405: out <= 16'hFEAD;    16'd45406: out <= 16'h0393;    16'd45407: out <= 16'h07D5;
    16'd45408: out <= 16'h0019;    16'd45409: out <= 16'h0625;    16'd45410: out <= 16'h036C;    16'd45411: out <= 16'h0214;
    16'd45412: out <= 16'h0046;    16'd45413: out <= 16'h0478;    16'd45414: out <= 16'h0933;    16'd45415: out <= 16'h0485;
    16'd45416: out <= 16'hFC4E;    16'd45417: out <= 16'h00CF;    16'd45418: out <= 16'hFDAA;    16'd45419: out <= 16'hFF5D;
    16'd45420: out <= 16'hFE8F;    16'd45421: out <= 16'h044A;    16'd45422: out <= 16'h0B84;    16'd45423: out <= 16'h0590;
    16'd45424: out <= 16'h027D;    16'd45425: out <= 16'h09CB;    16'd45426: out <= 16'h078A;    16'd45427: out <= 16'h0181;
    16'd45428: out <= 16'hFBF4;    16'd45429: out <= 16'h0126;    16'd45430: out <= 16'h0205;    16'd45431: out <= 16'h0668;
    16'd45432: out <= 16'h056A;    16'd45433: out <= 16'h0191;    16'd45434: out <= 16'h0451;    16'd45435: out <= 16'h0844;
    16'd45436: out <= 16'h08CC;    16'd45437: out <= 16'h0805;    16'd45438: out <= 16'h0139;    16'd45439: out <= 16'h0696;
    16'd45440: out <= 16'h0005;    16'd45441: out <= 16'hFD31;    16'd45442: out <= 16'hFF5F;    16'd45443: out <= 16'h05F8;
    16'd45444: out <= 16'h00D0;    16'd45445: out <= 16'h066E;    16'd45446: out <= 16'h0539;    16'd45447: out <= 16'h0DDD;
    16'd45448: out <= 16'h0334;    16'd45449: out <= 16'h06F5;    16'd45450: out <= 16'hFF88;    16'd45451: out <= 16'h06AF;
    16'd45452: out <= 16'h05F4;    16'd45453: out <= 16'h04BC;    16'd45454: out <= 16'hFE75;    16'd45455: out <= 16'h027F;
    16'd45456: out <= 16'h0D3E;    16'd45457: out <= 16'h0073;    16'd45458: out <= 16'h02BE;    16'd45459: out <= 16'h0063;
    16'd45460: out <= 16'h05A0;    16'd45461: out <= 16'h04CA;    16'd45462: out <= 16'h04EE;    16'd45463: out <= 16'h022F;
    16'd45464: out <= 16'hFD3D;    16'd45465: out <= 16'h0411;    16'd45466: out <= 16'h035F;    16'd45467: out <= 16'h0A6B;
    16'd45468: out <= 16'h0868;    16'd45469: out <= 16'h064A;    16'd45470: out <= 16'h02D9;    16'd45471: out <= 16'hFFB7;
    16'd45472: out <= 16'h0921;    16'd45473: out <= 16'hFAE7;    16'd45474: out <= 16'h02E7;    16'd45475: out <= 16'hFE1F;
    16'd45476: out <= 16'h0630;    16'd45477: out <= 16'h05A0;    16'd45478: out <= 16'h043D;    16'd45479: out <= 16'h0225;
    16'd45480: out <= 16'h0251;    16'd45481: out <= 16'h0369;    16'd45482: out <= 16'h0696;    16'd45483: out <= 16'h055C;
    16'd45484: out <= 16'h0698;    16'd45485: out <= 16'h0A7E;    16'd45486: out <= 16'h071B;    16'd45487: out <= 16'hFEED;
    16'd45488: out <= 16'h04E0;    16'd45489: out <= 16'h08B6;    16'd45490: out <= 16'h0546;    16'd45491: out <= 16'h0334;
    16'd45492: out <= 16'hFD9E;    16'd45493: out <= 16'h048D;    16'd45494: out <= 16'h0297;    16'd45495: out <= 16'h03DF;
    16'd45496: out <= 16'h0800;    16'd45497: out <= 16'h04B2;    16'd45498: out <= 16'h0753;    16'd45499: out <= 16'h00B5;
    16'd45500: out <= 16'h05FE;    16'd45501: out <= 16'hFE4D;    16'd45502: out <= 16'h0039;    16'd45503: out <= 16'h03DC;
    16'd45504: out <= 16'hFD36;    16'd45505: out <= 16'h0394;    16'd45506: out <= 16'h01C8;    16'd45507: out <= 16'h07BD;
    16'd45508: out <= 16'h0698;    16'd45509: out <= 16'h078D;    16'd45510: out <= 16'h08E4;    16'd45511: out <= 16'h07D2;
    16'd45512: out <= 16'h0563;    16'd45513: out <= 16'h096A;    16'd45514: out <= 16'h0198;    16'd45515: out <= 16'hFA97;
    16'd45516: out <= 16'h0311;    16'd45517: out <= 16'h0235;    16'd45518: out <= 16'hFFAD;    16'd45519: out <= 16'hFF01;
    16'd45520: out <= 16'hFA6A;    16'd45521: out <= 16'hFF85;    16'd45522: out <= 16'h0493;    16'd45523: out <= 16'hFC3F;
    16'd45524: out <= 16'h0367;    16'd45525: out <= 16'h0158;    16'd45526: out <= 16'h0000;    16'd45527: out <= 16'h025C;
    16'd45528: out <= 16'h0091;    16'd45529: out <= 16'h018A;    16'd45530: out <= 16'h006F;    16'd45531: out <= 16'h0296;
    16'd45532: out <= 16'hFF02;    16'd45533: out <= 16'h0186;    16'd45534: out <= 16'h04D6;    16'd45535: out <= 16'h0776;
    16'd45536: out <= 16'hFED2;    16'd45537: out <= 16'hF4E1;    16'd45538: out <= 16'hFD88;    16'd45539: out <= 16'h00B9;
    16'd45540: out <= 16'hFDF1;    16'd45541: out <= 16'h0416;    16'd45542: out <= 16'h029F;    16'd45543: out <= 16'h0923;
    16'd45544: out <= 16'hFF3E;    16'd45545: out <= 16'hFEAF;    16'd45546: out <= 16'hF93B;    16'd45547: out <= 16'hFFE0;
    16'd45548: out <= 16'hFBFE;    16'd45549: out <= 16'hF9A7;    16'd45550: out <= 16'hFF7B;    16'd45551: out <= 16'hFEA1;
    16'd45552: out <= 16'h0178;    16'd45553: out <= 16'h0264;    16'd45554: out <= 16'hFD26;    16'd45555: out <= 16'hFD4B;
    16'd45556: out <= 16'h054D;    16'd45557: out <= 16'hFCE8;    16'd45558: out <= 16'h0055;    16'd45559: out <= 16'h034F;
    16'd45560: out <= 16'h06DD;    16'd45561: out <= 16'h05FF;    16'd45562: out <= 16'h00A1;    16'd45563: out <= 16'h0184;
    16'd45564: out <= 16'hFADA;    16'd45565: out <= 16'hFD89;    16'd45566: out <= 16'h0943;    16'd45567: out <= 16'h00B4;
    16'd45568: out <= 16'hFBBE;    16'd45569: out <= 16'hFE1F;    16'd45570: out <= 16'hFA5E;    16'd45571: out <= 16'hFC4F;
    16'd45572: out <= 16'h0769;    16'd45573: out <= 16'h02A3;    16'd45574: out <= 16'h0126;    16'd45575: out <= 16'h007D;
    16'd45576: out <= 16'hFEB9;    16'd45577: out <= 16'h01C0;    16'd45578: out <= 16'hFEB7;    16'd45579: out <= 16'hFE4F;
    16'd45580: out <= 16'hFE77;    16'd45581: out <= 16'hFE88;    16'd45582: out <= 16'hFA1A;    16'd45583: out <= 16'hFF06;
    16'd45584: out <= 16'h0268;    16'd45585: out <= 16'h01AF;    16'd45586: out <= 16'h04DD;    16'd45587: out <= 16'h01D6;
    16'd45588: out <= 16'hFE1A;    16'd45589: out <= 16'hFFF1;    16'd45590: out <= 16'hFE8C;    16'd45591: out <= 16'hFF97;
    16'd45592: out <= 16'h0152;    16'd45593: out <= 16'h03D2;    16'd45594: out <= 16'h03E1;    16'd45595: out <= 16'hFFC3;
    16'd45596: out <= 16'hFDF1;    16'd45597: out <= 16'h016E;    16'd45598: out <= 16'h0247;    16'd45599: out <= 16'hFC31;
    16'd45600: out <= 16'hFD34;    16'd45601: out <= 16'h0508;    16'd45602: out <= 16'hFE3B;    16'd45603: out <= 16'hF9A2;
    16'd45604: out <= 16'h03B3;    16'd45605: out <= 16'h02E0;    16'd45606: out <= 16'h0798;    16'd45607: out <= 16'h0DCF;
    16'd45608: out <= 16'h002C;    16'd45609: out <= 16'h08D4;    16'd45610: out <= 16'h0150;    16'd45611: out <= 16'h02C7;
    16'd45612: out <= 16'h028A;    16'd45613: out <= 16'h057C;    16'd45614: out <= 16'h0510;    16'd45615: out <= 16'hFE93;
    16'd45616: out <= 16'hFFD8;    16'd45617: out <= 16'h019E;    16'd45618: out <= 16'h0152;    16'd45619: out <= 16'hFFB3;
    16'd45620: out <= 16'h09EE;    16'd45621: out <= 16'hFFA5;    16'd45622: out <= 16'h0493;    16'd45623: out <= 16'h0868;
    16'd45624: out <= 16'hFDCD;    16'd45625: out <= 16'h05EA;    16'd45626: out <= 16'h050A;    16'd45627: out <= 16'hFF36;
    16'd45628: out <= 16'hFEAB;    16'd45629: out <= 16'h0466;    16'd45630: out <= 16'h0577;    16'd45631: out <= 16'hFEC8;
    16'd45632: out <= 16'h03B4;    16'd45633: out <= 16'h04D3;    16'd45634: out <= 16'hFD2B;    16'd45635: out <= 16'h041C;
    16'd45636: out <= 16'h0729;    16'd45637: out <= 16'hFE25;    16'd45638: out <= 16'h0295;    16'd45639: out <= 16'h0BF4;
    16'd45640: out <= 16'h0304;    16'd45641: out <= 16'h065E;    16'd45642: out <= 16'h09A7;    16'd45643: out <= 16'h05D8;
    16'd45644: out <= 16'hFC71;    16'd45645: out <= 16'h0119;    16'd45646: out <= 16'hFBAE;    16'd45647: out <= 16'h047A;
    16'd45648: out <= 16'hFDD6;    16'd45649: out <= 16'h02B3;    16'd45650: out <= 16'h057E;    16'd45651: out <= 16'h0524;
    16'd45652: out <= 16'hFF55;    16'd45653: out <= 16'hFFEE;    16'd45654: out <= 16'h04D8;    16'd45655: out <= 16'h072F;
    16'd45656: out <= 16'h082E;    16'd45657: out <= 16'hFF23;    16'd45658: out <= 16'h07A5;    16'd45659: out <= 16'h041A;
    16'd45660: out <= 16'h0179;    16'd45661: out <= 16'h05CB;    16'd45662: out <= 16'h004B;    16'd45663: out <= 16'h0ABA;
    16'd45664: out <= 16'h02FE;    16'd45665: out <= 16'h0308;    16'd45666: out <= 16'h02E8;    16'd45667: out <= 16'h0C0F;
    16'd45668: out <= 16'h041E;    16'd45669: out <= 16'h04DC;    16'd45670: out <= 16'h03F2;    16'd45671: out <= 16'hFA3E;
    16'd45672: out <= 16'hFD9C;    16'd45673: out <= 16'h07AE;    16'd45674: out <= 16'h029F;    16'd45675: out <= 16'h0630;
    16'd45676: out <= 16'hF9BD;    16'd45677: out <= 16'h03FC;    16'd45678: out <= 16'hFB53;    16'd45679: out <= 16'hFE95;
    16'd45680: out <= 16'hFC54;    16'd45681: out <= 16'h0488;    16'd45682: out <= 16'h096D;    16'd45683: out <= 16'hFC40;
    16'd45684: out <= 16'h02AC;    16'd45685: out <= 16'h05AF;    16'd45686: out <= 16'hFEE3;    16'd45687: out <= 16'h0993;
    16'd45688: out <= 16'h043C;    16'd45689: out <= 16'hFE70;    16'd45690: out <= 16'h0BA1;    16'd45691: out <= 16'h09CD;
    16'd45692: out <= 16'h03E9;    16'd45693: out <= 16'hFE4B;    16'd45694: out <= 16'h092E;    16'd45695: out <= 16'h04D9;
    16'd45696: out <= 16'h07D1;    16'd45697: out <= 16'h0209;    16'd45698: out <= 16'h01C3;    16'd45699: out <= 16'h04C0;
    16'd45700: out <= 16'h0349;    16'd45701: out <= 16'h06F2;    16'd45702: out <= 16'h0670;    16'd45703: out <= 16'h00DB;
    16'd45704: out <= 16'h046F;    16'd45705: out <= 16'hFFF8;    16'd45706: out <= 16'h09CF;    16'd45707: out <= 16'h018F;
    16'd45708: out <= 16'h0809;    16'd45709: out <= 16'h0A3C;    16'd45710: out <= 16'h0180;    16'd45711: out <= 16'h0D10;
    16'd45712: out <= 16'h0846;    16'd45713: out <= 16'h07F5;    16'd45714: out <= 16'h0431;    16'd45715: out <= 16'h015D;
    16'd45716: out <= 16'h03C9;    16'd45717: out <= 16'h06FA;    16'd45718: out <= 16'h0342;    16'd45719: out <= 16'h079E;
    16'd45720: out <= 16'h0128;    16'd45721: out <= 16'hFD93;    16'd45722: out <= 16'hFAF3;    16'd45723: out <= 16'h06F3;
    16'd45724: out <= 16'h03DA;    16'd45725: out <= 16'h02F6;    16'd45726: out <= 16'h02DD;    16'd45727: out <= 16'h046C;
    16'd45728: out <= 16'h008F;    16'd45729: out <= 16'h027B;    16'd45730: out <= 16'hFE7B;    16'd45731: out <= 16'h0271;
    16'd45732: out <= 16'h084D;    16'd45733: out <= 16'h0538;    16'd45734: out <= 16'hFE4D;    16'd45735: out <= 16'h0874;
    16'd45736: out <= 16'h0614;    16'd45737: out <= 16'h0EC8;    16'd45738: out <= 16'hFE25;    16'd45739: out <= 16'hFD83;
    16'd45740: out <= 16'h05A5;    16'd45741: out <= 16'h0281;    16'd45742: out <= 16'hFC1E;    16'd45743: out <= 16'h0002;
    16'd45744: out <= 16'h0464;    16'd45745: out <= 16'h08BE;    16'd45746: out <= 16'h02F8;    16'd45747: out <= 16'h0A44;
    16'd45748: out <= 16'h0565;    16'd45749: out <= 16'h0AA7;    16'd45750: out <= 16'h019C;    16'd45751: out <= 16'h0511;
    16'd45752: out <= 16'h021B;    16'd45753: out <= 16'h0982;    16'd45754: out <= 16'hFFBA;    16'd45755: out <= 16'h0853;
    16'd45756: out <= 16'h045F;    16'd45757: out <= 16'h050F;    16'd45758: out <= 16'h0A25;    16'd45759: out <= 16'h01F6;
    16'd45760: out <= 16'h0574;    16'd45761: out <= 16'h0020;    16'd45762: out <= 16'h0069;    16'd45763: out <= 16'h094C;
    16'd45764: out <= 16'h01F7;    16'd45765: out <= 16'hF998;    16'd45766: out <= 16'h0530;    16'd45767: out <= 16'h048E;
    16'd45768: out <= 16'h09FA;    16'd45769: out <= 16'h0431;    16'd45770: out <= 16'h09AF;    16'd45771: out <= 16'hFB4D;
    16'd45772: out <= 16'hFEF7;    16'd45773: out <= 16'hF777;    16'd45774: out <= 16'hFC59;    16'd45775: out <= 16'h04FC;
    16'd45776: out <= 16'hF7C0;    16'd45777: out <= 16'hFEE1;    16'd45778: out <= 16'h02F5;    16'd45779: out <= 16'hF8AB;
    16'd45780: out <= 16'h0198;    16'd45781: out <= 16'hFBCE;    16'd45782: out <= 16'hF872;    16'd45783: out <= 16'h025E;
    16'd45784: out <= 16'h02BC;    16'd45785: out <= 16'h0131;    16'd45786: out <= 16'hF981;    16'd45787: out <= 16'hFB70;
    16'd45788: out <= 16'h00EC;    16'd45789: out <= 16'h0003;    16'd45790: out <= 16'h0105;    16'd45791: out <= 16'h0227;
    16'd45792: out <= 16'hFE78;    16'd45793: out <= 16'hFFEC;    16'd45794: out <= 16'hF98E;    16'd45795: out <= 16'hFFC0;
    16'd45796: out <= 16'hFED4;    16'd45797: out <= 16'h0292;    16'd45798: out <= 16'hFEC6;    16'd45799: out <= 16'hFD46;
    16'd45800: out <= 16'h04DE;    16'd45801: out <= 16'h0954;    16'd45802: out <= 16'h04B8;    16'd45803: out <= 16'hF9B9;
    16'd45804: out <= 16'hFAC7;    16'd45805: out <= 16'hFE1A;    16'd45806: out <= 16'h01C3;    16'd45807: out <= 16'hF812;
    16'd45808: out <= 16'h0056;    16'd45809: out <= 16'h000A;    16'd45810: out <= 16'h0385;    16'd45811: out <= 16'h02DF;
    16'd45812: out <= 16'hF96D;    16'd45813: out <= 16'h03A1;    16'd45814: out <= 16'h0468;    16'd45815: out <= 16'hFA3F;
    16'd45816: out <= 16'hFA22;    16'd45817: out <= 16'h0667;    16'd45818: out <= 16'hFA3A;    16'd45819: out <= 16'h0454;
    16'd45820: out <= 16'h02C7;    16'd45821: out <= 16'h05A4;    16'd45822: out <= 16'h0636;    16'd45823: out <= 16'h008E;
    16'd45824: out <= 16'h01CF;    16'd45825: out <= 16'h017C;    16'd45826: out <= 16'h01C4;    16'd45827: out <= 16'hFF27;
    16'd45828: out <= 16'hFD7C;    16'd45829: out <= 16'h01D6;    16'd45830: out <= 16'h0081;    16'd45831: out <= 16'h03F4;
    16'd45832: out <= 16'hFDAE;    16'd45833: out <= 16'h01C3;    16'd45834: out <= 16'hF853;    16'd45835: out <= 16'h0068;
    16'd45836: out <= 16'hFD66;    16'd45837: out <= 16'h0196;    16'd45838: out <= 16'hFBEA;    16'd45839: out <= 16'h002F;
    16'd45840: out <= 16'h019C;    16'd45841: out <= 16'hFE1E;    16'd45842: out <= 16'h03E9;    16'd45843: out <= 16'hFF18;
    16'd45844: out <= 16'hFDF7;    16'd45845: out <= 16'hF98E;    16'd45846: out <= 16'hFFA1;    16'd45847: out <= 16'h0302;
    16'd45848: out <= 16'h042F;    16'd45849: out <= 16'h00B4;    16'd45850: out <= 16'hFA47;    16'd45851: out <= 16'h0316;
    16'd45852: out <= 16'h0493;    16'd45853: out <= 16'hFE1E;    16'd45854: out <= 16'h0231;    16'd45855: out <= 16'hFF0B;
    16'd45856: out <= 16'hFE4E;    16'd45857: out <= 16'h06E0;    16'd45858: out <= 16'h00A4;    16'd45859: out <= 16'h0434;
    16'd45860: out <= 16'h02BF;    16'd45861: out <= 16'h0097;    16'd45862: out <= 16'h05B0;    16'd45863: out <= 16'h00BC;
    16'd45864: out <= 16'hFFC5;    16'd45865: out <= 16'h05FF;    16'd45866: out <= 16'h02A3;    16'd45867: out <= 16'h032B;
    16'd45868: out <= 16'h059C;    16'd45869: out <= 16'h0487;    16'd45870: out <= 16'h027E;    16'd45871: out <= 16'h014D;
    16'd45872: out <= 16'h03AB;    16'd45873: out <= 16'h0859;    16'd45874: out <= 16'hFF04;    16'd45875: out <= 16'h0478;
    16'd45876: out <= 16'h0951;    16'd45877: out <= 16'h0395;    16'd45878: out <= 16'h075D;    16'd45879: out <= 16'h071E;
    16'd45880: out <= 16'h076A;    16'd45881: out <= 16'h06D2;    16'd45882: out <= 16'h07ED;    16'd45883: out <= 16'h0618;
    16'd45884: out <= 16'h0270;    16'd45885: out <= 16'h0902;    16'd45886: out <= 16'h061C;    16'd45887: out <= 16'h03E5;
    16'd45888: out <= 16'hFF23;    16'd45889: out <= 16'h0500;    16'd45890: out <= 16'h0858;    16'd45891: out <= 16'h0CB8;
    16'd45892: out <= 16'h0C41;    16'd45893: out <= 16'h0179;    16'd45894: out <= 16'h0556;    16'd45895: out <= 16'h02A6;
    16'd45896: out <= 16'h0413;    16'd45897: out <= 16'h0370;    16'd45898: out <= 16'hFECF;    16'd45899: out <= 16'h010E;
    16'd45900: out <= 16'hFD83;    16'd45901: out <= 16'h0228;    16'd45902: out <= 16'hFBC7;    16'd45903: out <= 16'h028A;
    16'd45904: out <= 16'h0118;    16'd45905: out <= 16'h00CB;    16'd45906: out <= 16'h02ED;    16'd45907: out <= 16'h0099;
    16'd45908: out <= 16'hF94A;    16'd45909: out <= 16'h075B;    16'd45910: out <= 16'hFE87;    16'd45911: out <= 16'h0094;
    16'd45912: out <= 16'h00D6;    16'd45913: out <= 16'h06E4;    16'd45914: out <= 16'h0508;    16'd45915: out <= 16'h0679;
    16'd45916: out <= 16'h0933;    16'd45917: out <= 16'h0BC5;    16'd45918: out <= 16'h065A;    16'd45919: out <= 16'h0756;
    16'd45920: out <= 16'h032D;    16'd45921: out <= 16'h069F;    16'd45922: out <= 16'hFFAB;    16'd45923: out <= 16'h0273;
    16'd45924: out <= 16'h0045;    16'd45925: out <= 16'hFF23;    16'd45926: out <= 16'hFEAC;    16'd45927: out <= 16'hF6BF;
    16'd45928: out <= 16'hFBEF;    16'd45929: out <= 16'h0488;    16'd45930: out <= 16'h073D;    16'd45931: out <= 16'hFFF9;
    16'd45932: out <= 16'h002C;    16'd45933: out <= 16'h0178;    16'd45934: out <= 16'h029E;    16'd45935: out <= 16'hF99A;
    16'd45936: out <= 16'h023A;    16'd45937: out <= 16'h004D;    16'd45938: out <= 16'h0592;    16'd45939: out <= 16'hFEDA;
    16'd45940: out <= 16'hFE33;    16'd45941: out <= 16'h00DF;    16'd45942: out <= 16'hFD91;    16'd45943: out <= 16'h0629;
    16'd45944: out <= 16'h0588;    16'd45945: out <= 16'hF9E1;    16'd45946: out <= 16'hFD5D;    16'd45947: out <= 16'hFF8F;
    16'd45948: out <= 16'h004F;    16'd45949: out <= 16'h00C4;    16'd45950: out <= 16'h0016;    16'd45951: out <= 16'h0074;
    16'd45952: out <= 16'hFCE2;    16'd45953: out <= 16'h0C73;    16'd45954: out <= 16'h0651;    16'd45955: out <= 16'h0658;
    16'd45956: out <= 16'h033B;    16'd45957: out <= 16'h08CF;    16'd45958: out <= 16'h082A;    16'd45959: out <= 16'h07D8;
    16'd45960: out <= 16'h0409;    16'd45961: out <= 16'h010A;    16'd45962: out <= 16'h0259;    16'd45963: out <= 16'h02C5;
    16'd45964: out <= 16'h09C6;    16'd45965: out <= 16'hFAB4;    16'd45966: out <= 16'h05A3;    16'd45967: out <= 16'h044B;
    16'd45968: out <= 16'h01BA;    16'd45969: out <= 16'h0522;    16'd45970: out <= 16'h053A;    16'd45971: out <= 16'h04E5;
    16'd45972: out <= 16'h0627;    16'd45973: out <= 16'h0109;    16'd45974: out <= 16'h0E83;    16'd45975: out <= 16'h03D3;
    16'd45976: out <= 16'h027A;    16'd45977: out <= 16'h057F;    16'd45978: out <= 16'h0952;    16'd45979: out <= 16'h02B7;
    16'd45980: out <= 16'h07D6;    16'd45981: out <= 16'hFEED;    16'd45982: out <= 16'h08A0;    16'd45983: out <= 16'hFE74;
    16'd45984: out <= 16'hFA32;    16'd45985: out <= 16'h0966;    16'd45986: out <= 16'h05B0;    16'd45987: out <= 16'h06E0;
    16'd45988: out <= 16'hFF92;    16'd45989: out <= 16'h0387;    16'd45990: out <= 16'h060C;    16'd45991: out <= 16'hFE26;
    16'd45992: out <= 16'h0762;    16'd45993: out <= 16'h0BCD;    16'd45994: out <= 16'hFFE8;    16'd45995: out <= 16'h07B7;
    16'd45996: out <= 16'h0230;    16'd45997: out <= 16'h0883;    16'd45998: out <= 16'h00FD;    16'd45999: out <= 16'h0920;
    16'd46000: out <= 16'h0839;    16'd46001: out <= 16'h0427;    16'd46002: out <= 16'h04C0;    16'd46003: out <= 16'h040F;
    16'd46004: out <= 16'h0461;    16'd46005: out <= 16'hFBF0;    16'd46006: out <= 16'h0380;    16'd46007: out <= 16'h00A4;
    16'd46008: out <= 16'h0376;    16'd46009: out <= 16'hFE6A;    16'd46010: out <= 16'hFEFE;    16'd46011: out <= 16'hFBB1;
    16'd46012: out <= 16'h0033;    16'd46013: out <= 16'h0999;    16'd46014: out <= 16'h074B;    16'd46015: out <= 16'h06B5;
    16'd46016: out <= 16'h03D5;    16'd46017: out <= 16'hFE0C;    16'd46018: out <= 16'h0012;    16'd46019: out <= 16'h061D;
    16'd46020: out <= 16'h04D2;    16'd46021: out <= 16'h0131;    16'd46022: out <= 16'h072E;    16'd46023: out <= 16'hFCDD;
    16'd46024: out <= 16'h04CA;    16'd46025: out <= 16'h0510;    16'd46026: out <= 16'h03DD;    16'd46027: out <= 16'h02EB;
    16'd46028: out <= 16'hFDA5;    16'd46029: out <= 16'h00CF;    16'd46030: out <= 16'hFE25;    16'd46031: out <= 16'hFCA0;
    16'd46032: out <= 16'hFFB8;    16'd46033: out <= 16'h0085;    16'd46034: out <= 16'hFDC7;    16'd46035: out <= 16'hFE59;
    16'd46036: out <= 16'h020F;    16'd46037: out <= 16'hFB6D;    16'd46038: out <= 16'hFD4A;    16'd46039: out <= 16'hFE2B;
    16'd46040: out <= 16'hFC88;    16'd46041: out <= 16'hFC9D;    16'd46042: out <= 16'hFF07;    16'd46043: out <= 16'h01C9;
    16'd46044: out <= 16'hFDAD;    16'd46045: out <= 16'h034C;    16'd46046: out <= 16'h0253;    16'd46047: out <= 16'h0955;
    16'd46048: out <= 16'hFD90;    16'd46049: out <= 16'h0138;    16'd46050: out <= 16'h0539;    16'd46051: out <= 16'hFA4F;
    16'd46052: out <= 16'hF984;    16'd46053: out <= 16'hFEAF;    16'd46054: out <= 16'h00E0;    16'd46055: out <= 16'h067E;
    16'd46056: out <= 16'h05A1;    16'd46057: out <= 16'hFF13;    16'd46058: out <= 16'h0022;    16'd46059: out <= 16'h00EC;
    16'd46060: out <= 16'h0178;    16'd46061: out <= 16'h0074;    16'd46062: out <= 16'h013F;    16'd46063: out <= 16'hFE1E;
    16'd46064: out <= 16'hFA66;    16'd46065: out <= 16'h02D3;    16'd46066: out <= 16'h029B;    16'd46067: out <= 16'hFDFF;
    16'd46068: out <= 16'hFF2C;    16'd46069: out <= 16'h0469;    16'd46070: out <= 16'hFABE;    16'd46071: out <= 16'h004E;
    16'd46072: out <= 16'hFCC6;    16'd46073: out <= 16'hFE21;    16'd46074: out <= 16'hFE82;    16'd46075: out <= 16'h0064;
    16'd46076: out <= 16'hFF95;    16'd46077: out <= 16'h0053;    16'd46078: out <= 16'hFE6C;    16'd46079: out <= 16'hFF8D;
    16'd46080: out <= 16'h0438;    16'd46081: out <= 16'h009E;    16'd46082: out <= 16'h00FF;    16'd46083: out <= 16'hFC59;
    16'd46084: out <= 16'h001A;    16'd46085: out <= 16'hFDD4;    16'd46086: out <= 16'hFE04;    16'd46087: out <= 16'h01A2;
    16'd46088: out <= 16'h0248;    16'd46089: out <= 16'hFCC5;    16'd46090: out <= 16'h0175;    16'd46091: out <= 16'hFEF9;
    16'd46092: out <= 16'hFAFC;    16'd46093: out <= 16'hFD8E;    16'd46094: out <= 16'hFE7B;    16'd46095: out <= 16'h023D;
    16'd46096: out <= 16'h0192;    16'd46097: out <= 16'hFDFB;    16'd46098: out <= 16'h062A;    16'd46099: out <= 16'hFBA2;
    16'd46100: out <= 16'h02D4;    16'd46101: out <= 16'h013C;    16'd46102: out <= 16'hFEBE;    16'd46103: out <= 16'h060E;
    16'd46104: out <= 16'h0129;    16'd46105: out <= 16'h02BD;    16'd46106: out <= 16'h025F;    16'd46107: out <= 16'h016C;
    16'd46108: out <= 16'h0274;    16'd46109: out <= 16'h007E;    16'd46110: out <= 16'h0645;    16'd46111: out <= 16'h004C;
    16'd46112: out <= 16'hFE17;    16'd46113: out <= 16'hFC3C;    16'd46114: out <= 16'h039B;    16'd46115: out <= 16'hFC48;
    16'd46116: out <= 16'hFD09;    16'd46117: out <= 16'h06CF;    16'd46118: out <= 16'h0729;    16'd46119: out <= 16'h0A77;
    16'd46120: out <= 16'hFFE2;    16'd46121: out <= 16'hFDA7;    16'd46122: out <= 16'h04FE;    16'd46123: out <= 16'h0940;
    16'd46124: out <= 16'hFFD6;    16'd46125: out <= 16'h0503;    16'd46126: out <= 16'h06A4;    16'd46127: out <= 16'h0E0E;
    16'd46128: out <= 16'h04B4;    16'd46129: out <= 16'h055E;    16'd46130: out <= 16'h04B7;    16'd46131: out <= 16'hFBD0;
    16'd46132: out <= 16'h0245;    16'd46133: out <= 16'h017B;    16'd46134: out <= 16'h0221;    16'd46135: out <= 16'h0154;
    16'd46136: out <= 16'h0814;    16'd46137: out <= 16'h055D;    16'd46138: out <= 16'h05E9;    16'd46139: out <= 16'h0381;
    16'd46140: out <= 16'hFFCC;    16'd46141: out <= 16'h024C;    16'd46142: out <= 16'h0457;    16'd46143: out <= 16'h02FF;
    16'd46144: out <= 16'h02BE;    16'd46145: out <= 16'h006D;    16'd46146: out <= 16'h07DA;    16'd46147: out <= 16'h01BD;
    16'd46148: out <= 16'h0103;    16'd46149: out <= 16'h047D;    16'd46150: out <= 16'h005B;    16'd46151: out <= 16'h053F;
    16'd46152: out <= 16'hFF86;    16'd46153: out <= 16'h01C7;    16'd46154: out <= 16'h021A;    16'd46155: out <= 16'h0195;
    16'd46156: out <= 16'h024D;    16'd46157: out <= 16'h0314;    16'd46158: out <= 16'hFD22;    16'd46159: out <= 16'h0010;
    16'd46160: out <= 16'h02FA;    16'd46161: out <= 16'hFEA2;    16'd46162: out <= 16'hFED4;    16'd46163: out <= 16'h0015;
    16'd46164: out <= 16'h03ED;    16'd46165: out <= 16'h04AC;    16'd46166: out <= 16'h0478;    16'd46167: out <= 16'hFC60;
    16'd46168: out <= 16'hFF9F;    16'd46169: out <= 16'hFD48;    16'd46170: out <= 16'h0052;    16'd46171: out <= 16'hFFF4;
    16'd46172: out <= 16'h0078;    16'd46173: out <= 16'h061D;    16'd46174: out <= 16'hFF7E;    16'd46175: out <= 16'hFFA1;
    16'd46176: out <= 16'h001D;    16'd46177: out <= 16'h09EC;    16'd46178: out <= 16'h0185;    16'd46179: out <= 16'h081A;
    16'd46180: out <= 16'h06DE;    16'd46181: out <= 16'hFE4F;    16'd46182: out <= 16'h0444;    16'd46183: out <= 16'h0083;
    16'd46184: out <= 16'hFC65;    16'd46185: out <= 16'h042E;    16'd46186: out <= 16'h044A;    16'd46187: out <= 16'hFC68;
    16'd46188: out <= 16'hF965;    16'd46189: out <= 16'h05D8;    16'd46190: out <= 16'hFAD8;    16'd46191: out <= 16'h0108;
    16'd46192: out <= 16'hFD09;    16'd46193: out <= 16'h01F2;    16'd46194: out <= 16'hFF0A;    16'd46195: out <= 16'hFD86;
    16'd46196: out <= 16'hFA00;    16'd46197: out <= 16'hFE66;    16'd46198: out <= 16'h004C;    16'd46199: out <= 16'hFB4B;
    16'd46200: out <= 16'hF9F4;    16'd46201: out <= 16'h0085;    16'd46202: out <= 16'hFC63;    16'd46203: out <= 16'h02EC;
    16'd46204: out <= 16'hFE44;    16'd46205: out <= 16'h0560;    16'd46206: out <= 16'h0170;    16'd46207: out <= 16'hFFE7;
    16'd46208: out <= 16'h00D3;    16'd46209: out <= 16'h02B6;    16'd46210: out <= 16'h05B9;    16'd46211: out <= 16'hFFE5;
    16'd46212: out <= 16'h0007;    16'd46213: out <= 16'h06E7;    16'd46214: out <= 16'h0757;    16'd46215: out <= 16'h010B;
    16'd46216: out <= 16'h029E;    16'd46217: out <= 16'h058A;    16'd46218: out <= 16'h0379;    16'd46219: out <= 16'h0001;
    16'd46220: out <= 16'h003A;    16'd46221: out <= 16'h0122;    16'd46222: out <= 16'hFEDC;    16'd46223: out <= 16'h0353;
    16'd46224: out <= 16'h08C8;    16'd46225: out <= 16'hFC67;    16'd46226: out <= 16'hFFF6;    16'd46227: out <= 16'h0143;
    16'd46228: out <= 16'h054D;    16'd46229: out <= 16'hFD47;    16'd46230: out <= 16'h096B;    16'd46231: out <= 16'hFE3E;
    16'd46232: out <= 16'h0671;    16'd46233: out <= 16'h0A90;    16'd46234: out <= 16'h0A24;    16'd46235: out <= 16'h0278;
    16'd46236: out <= 16'h049A;    16'd46237: out <= 16'h02E7;    16'd46238: out <= 16'h0460;    16'd46239: out <= 16'h07EB;
    16'd46240: out <= 16'h063A;    16'd46241: out <= 16'h006A;    16'd46242: out <= 16'h05B9;    16'd46243: out <= 16'h0889;
    16'd46244: out <= 16'h0446;    16'd46245: out <= 16'h0533;    16'd46246: out <= 16'h0940;    16'd46247: out <= 16'h0350;
    16'd46248: out <= 16'h0608;    16'd46249: out <= 16'h05A1;    16'd46250: out <= 16'h035B;    16'd46251: out <= 16'hFE90;
    16'd46252: out <= 16'h093E;    16'd46253: out <= 16'h091C;    16'd46254: out <= 16'hFC86;    16'd46255: out <= 16'h08D8;
    16'd46256: out <= 16'h0530;    16'd46257: out <= 16'h07B8;    16'd46258: out <= 16'hFFEA;    16'd46259: out <= 16'h0634;
    16'd46260: out <= 16'h0931;    16'd46261: out <= 16'h073D;    16'd46262: out <= 16'h0330;    16'd46263: out <= 16'h0668;
    16'd46264: out <= 16'hFE94;    16'd46265: out <= 16'hFCA7;    16'd46266: out <= 16'h0232;    16'd46267: out <= 16'h051E;
    16'd46268: out <= 16'h02E8;    16'd46269: out <= 16'hFEBB;    16'd46270: out <= 16'h0873;    16'd46271: out <= 16'h024B;
    16'd46272: out <= 16'h04E9;    16'd46273: out <= 16'h01A0;    16'd46274: out <= 16'h0208;    16'd46275: out <= 16'h04BD;
    16'd46276: out <= 16'hFEDD;    16'd46277: out <= 16'h017E;    16'd46278: out <= 16'h04A2;    16'd46279: out <= 16'h05E4;
    16'd46280: out <= 16'h0617;    16'd46281: out <= 16'h0112;    16'd46282: out <= 16'h006D;    16'd46283: out <= 16'hFBC7;
    16'd46284: out <= 16'h0BAB;    16'd46285: out <= 16'hFE9C;    16'd46286: out <= 16'hFD3B;    16'd46287: out <= 16'h04C5;
    16'd46288: out <= 16'hFF66;    16'd46289: out <= 16'hFF35;    16'd46290: out <= 16'hFEC0;    16'd46291: out <= 16'h0087;
    16'd46292: out <= 16'hFC23;    16'd46293: out <= 16'h0394;    16'd46294: out <= 16'h0228;    16'd46295: out <= 16'h057F;
    16'd46296: out <= 16'hFBD6;    16'd46297: out <= 16'h02D2;    16'd46298: out <= 16'hFE6C;    16'd46299: out <= 16'hFFE8;
    16'd46300: out <= 16'hFF2A;    16'd46301: out <= 16'h0540;    16'd46302: out <= 16'h01B0;    16'd46303: out <= 16'h008D;
    16'd46304: out <= 16'h041A;    16'd46305: out <= 16'h000B;    16'd46306: out <= 16'h0792;    16'd46307: out <= 16'hF9CC;
    16'd46308: out <= 16'h0041;    16'd46309: out <= 16'hFCCD;    16'd46310: out <= 16'hFA04;    16'd46311: out <= 16'h0498;
    16'd46312: out <= 16'h04FD;    16'd46313: out <= 16'h074D;    16'd46314: out <= 16'h029F;    16'd46315: out <= 16'h05B9;
    16'd46316: out <= 16'h0155;    16'd46317: out <= 16'h0A04;    16'd46318: out <= 16'h0420;    16'd46319: out <= 16'hFFB8;
    16'd46320: out <= 16'h010B;    16'd46321: out <= 16'hFA50;    16'd46322: out <= 16'h038B;    16'd46323: out <= 16'h001A;
    16'd46324: out <= 16'h0195;    16'd46325: out <= 16'h06A7;    16'd46326: out <= 16'hFF9A;    16'd46327: out <= 16'hFD11;
    16'd46328: out <= 16'hFE32;    16'd46329: out <= 16'hFC43;    16'd46330: out <= 16'h00B8;    16'd46331: out <= 16'h02DE;
    16'd46332: out <= 16'hF9EA;    16'd46333: out <= 16'h0731;    16'd46334: out <= 16'h008D;    16'd46335: out <= 16'hFF81;
    16'd46336: out <= 16'hFC84;    16'd46337: out <= 16'hFBCC;    16'd46338: out <= 16'h019A;    16'd46339: out <= 16'hFF00;
    16'd46340: out <= 16'h0122;    16'd46341: out <= 16'h0289;    16'd46342: out <= 16'h0494;    16'd46343: out <= 16'hFCE5;
    16'd46344: out <= 16'hFB99;    16'd46345: out <= 16'hFF1D;    16'd46346: out <= 16'h00D6;    16'd46347: out <= 16'h02CF;
    16'd46348: out <= 16'h0782;    16'd46349: out <= 16'h05B0;    16'd46350: out <= 16'hFB5D;    16'd46351: out <= 16'hFD82;
    16'd46352: out <= 16'h0123;    16'd46353: out <= 16'hFF6D;    16'd46354: out <= 16'hFA2C;    16'd46355: out <= 16'h05D8;
    16'd46356: out <= 16'hFF7B;    16'd46357: out <= 16'h00B5;    16'd46358: out <= 16'h02D9;    16'd46359: out <= 16'hFF28;
    16'd46360: out <= 16'h00AC;    16'd46361: out <= 16'hFF47;    16'd46362: out <= 16'h0084;    16'd46363: out <= 16'hF9F7;
    16'd46364: out <= 16'hFFFA;    16'd46365: out <= 16'hFC68;    16'd46366: out <= 16'h054D;    16'd46367: out <= 16'h04C0;
    16'd46368: out <= 16'hFAA2;    16'd46369: out <= 16'h0608;    16'd46370: out <= 16'h022B;    16'd46371: out <= 16'hFCBD;
    16'd46372: out <= 16'hF505;    16'd46373: out <= 16'hFAFD;    16'd46374: out <= 16'h0345;    16'd46375: out <= 16'h0113;
    16'd46376: out <= 16'h07B0;    16'd46377: out <= 16'h037B;    16'd46378: out <= 16'hFD5B;    16'd46379: out <= 16'h005C;
    16'd46380: out <= 16'hFEA3;    16'd46381: out <= 16'h0500;    16'd46382: out <= 16'hF991;    16'd46383: out <= 16'hFF3D;
    16'd46384: out <= 16'h02B2;    16'd46385: out <= 16'hFFA2;    16'd46386: out <= 16'hF6BA;    16'd46387: out <= 16'h04FC;
    16'd46388: out <= 16'h058C;    16'd46389: out <= 16'h082D;    16'd46390: out <= 16'h0390;    16'd46391: out <= 16'h005D;
    16'd46392: out <= 16'h01A6;    16'd46393: out <= 16'h0C26;    16'd46394: out <= 16'h07C3;    16'd46395: out <= 16'h0095;
    16'd46396: out <= 16'h0A2C;    16'd46397: out <= 16'h0581;    16'd46398: out <= 16'h0598;    16'd46399: out <= 16'h005F;
    16'd46400: out <= 16'h0A44;    16'd46401: out <= 16'h022C;    16'd46402: out <= 16'h04C7;    16'd46403: out <= 16'h0408;
    16'd46404: out <= 16'h004B;    16'd46405: out <= 16'h03E2;    16'd46406: out <= 16'h021B;    16'd46407: out <= 16'h05AA;
    16'd46408: out <= 16'h06E6;    16'd46409: out <= 16'h01B4;    16'd46410: out <= 16'hFF13;    16'd46411: out <= 16'h0204;
    16'd46412: out <= 16'hFFBA;    16'd46413: out <= 16'h0008;    16'd46414: out <= 16'hFDE4;    16'd46415: out <= 16'hFB1C;
    16'd46416: out <= 16'hF955;    16'd46417: out <= 16'hF86E;    16'd46418: out <= 16'hFB2D;    16'd46419: out <= 16'hFD67;
    16'd46420: out <= 16'h0446;    16'd46421: out <= 16'hFC02;    16'd46422: out <= 16'h03E1;    16'd46423: out <= 16'h0526;
    16'd46424: out <= 16'hF990;    16'd46425: out <= 16'h0701;    16'd46426: out <= 16'h0357;    16'd46427: out <= 16'hFE2F;
    16'd46428: out <= 16'hFFF7;    16'd46429: out <= 16'hFE0B;    16'd46430: out <= 16'h00C9;    16'd46431: out <= 16'hFDD6;
    16'd46432: out <= 16'h03C0;    16'd46433: out <= 16'hFE07;    16'd46434: out <= 16'hFE94;    16'd46435: out <= 16'hFD64;
    16'd46436: out <= 16'hFF43;    16'd46437: out <= 16'h00B1;    16'd46438: out <= 16'hFFFB;    16'd46439: out <= 16'hFC58;
    16'd46440: out <= 16'hF828;    16'd46441: out <= 16'h0161;    16'd46442: out <= 16'h032F;    16'd46443: out <= 16'h00F3;
    16'd46444: out <= 16'hFE92;    16'd46445: out <= 16'hFCEF;    16'd46446: out <= 16'hFAFB;    16'd46447: out <= 16'hFD61;
    16'd46448: out <= 16'hFB05;    16'd46449: out <= 16'hFA45;    16'd46450: out <= 16'hFE2F;    16'd46451: out <= 16'h0A43;
    16'd46452: out <= 16'h0314;    16'd46453: out <= 16'h00E8;    16'd46454: out <= 16'hFC4B;    16'd46455: out <= 16'hFCB4;
    16'd46456: out <= 16'h017D;    16'd46457: out <= 16'hF9B4;    16'd46458: out <= 16'hFCBF;    16'd46459: out <= 16'hFED9;
    16'd46460: out <= 16'h006E;    16'd46461: out <= 16'hFCA2;    16'd46462: out <= 16'h0995;    16'd46463: out <= 16'h0141;
    16'd46464: out <= 16'hFF30;    16'd46465: out <= 16'h03B1;    16'd46466: out <= 16'h08BE;    16'd46467: out <= 16'hFE6F;
    16'd46468: out <= 16'hFE1B;    16'd46469: out <= 16'h0755;    16'd46470: out <= 16'h0DBE;    16'd46471: out <= 16'h0484;
    16'd46472: out <= 16'h0441;    16'd46473: out <= 16'h0567;    16'd46474: out <= 16'h047F;    16'd46475: out <= 16'h091E;
    16'd46476: out <= 16'h01FD;    16'd46477: out <= 16'h0DE5;    16'd46478: out <= 16'h03F8;    16'd46479: out <= 16'h0689;
    16'd46480: out <= 16'h0471;    16'd46481: out <= 16'h04F8;    16'd46482: out <= 16'h07E7;    16'd46483: out <= 16'hFF50;
    16'd46484: out <= 16'h028B;    16'd46485: out <= 16'h0ACA;    16'd46486: out <= 16'h04F4;    16'd46487: out <= 16'h02E8;
    16'd46488: out <= 16'hFDE1;    16'd46489: out <= 16'hFEB7;    16'd46490: out <= 16'h0A5B;    16'd46491: out <= 16'hFF4F;
    16'd46492: out <= 16'h0240;    16'd46493: out <= 16'hFE64;    16'd46494: out <= 16'h0585;    16'd46495: out <= 16'h0BD0;
    16'd46496: out <= 16'h0017;    16'd46497: out <= 16'h0350;    16'd46498: out <= 16'h0C04;    16'd46499: out <= 16'h0384;
    16'd46500: out <= 16'h0558;    16'd46501: out <= 16'h04F4;    16'd46502: out <= 16'h0026;    16'd46503: out <= 16'h061E;
    16'd46504: out <= 16'h0558;    16'd46505: out <= 16'h02A7;    16'd46506: out <= 16'hFDD1;    16'd46507: out <= 16'hFDA7;
    16'd46508: out <= 16'h0407;    16'd46509: out <= 16'h0709;    16'd46510: out <= 16'h0116;    16'd46511: out <= 16'h04F0;
    16'd46512: out <= 16'h063A;    16'd46513: out <= 16'h04B8;    16'd46514: out <= 16'h0485;    16'd46515: out <= 16'h0CCB;
    16'd46516: out <= 16'h0773;    16'd46517: out <= 16'h0483;    16'd46518: out <= 16'h008B;    16'd46519: out <= 16'h0090;
    16'd46520: out <= 16'h03A8;    16'd46521: out <= 16'h0201;    16'd46522: out <= 16'h0398;    16'd46523: out <= 16'hFC7C;
    16'd46524: out <= 16'hFD1B;    16'd46525: out <= 16'h05C1;    16'd46526: out <= 16'h060A;    16'd46527: out <= 16'h0174;
    16'd46528: out <= 16'h0503;    16'd46529: out <= 16'hFDB6;    16'd46530: out <= 16'h0079;    16'd46531: out <= 16'h0055;
    16'd46532: out <= 16'h0C54;    16'd46533: out <= 16'h05D5;    16'd46534: out <= 16'h05C0;    16'd46535: out <= 16'h0486;
    16'd46536: out <= 16'h02FE;    16'd46537: out <= 16'hFF3D;    16'd46538: out <= 16'h01F5;    16'd46539: out <= 16'h02EA;
    16'd46540: out <= 16'hFE86;    16'd46541: out <= 16'hF961;    16'd46542: out <= 16'h0592;    16'd46543: out <= 16'hFE17;
    16'd46544: out <= 16'h001D;    16'd46545: out <= 16'h0048;    16'd46546: out <= 16'h05A5;    16'd46547: out <= 16'hFE81;
    16'd46548: out <= 16'hFA44;    16'd46549: out <= 16'h01B2;    16'd46550: out <= 16'h0907;    16'd46551: out <= 16'h0040;
    16'd46552: out <= 16'h00E2;    16'd46553: out <= 16'hFE2A;    16'd46554: out <= 16'h0028;    16'd46555: out <= 16'hFE9D;
    16'd46556: out <= 16'h0572;    16'd46557: out <= 16'h0936;    16'd46558: out <= 16'h005F;    16'd46559: out <= 16'hFC86;
    16'd46560: out <= 16'hFFDB;    16'd46561: out <= 16'hFEC7;    16'd46562: out <= 16'h02AC;    16'd46563: out <= 16'h03AC;
    16'd46564: out <= 16'h0198;    16'd46565: out <= 16'hFFC0;    16'd46566: out <= 16'h07E1;    16'd46567: out <= 16'h0BA2;
    16'd46568: out <= 16'h032A;    16'd46569: out <= 16'hFBCF;    16'd46570: out <= 16'h0296;    16'd46571: out <= 16'hFA69;
    16'd46572: out <= 16'hF82C;    16'd46573: out <= 16'hFC2A;    16'd46574: out <= 16'hFD32;    16'd46575: out <= 16'h0365;
    16'd46576: out <= 16'hFA4C;    16'd46577: out <= 16'h01E7;    16'd46578: out <= 16'hFED9;    16'd46579: out <= 16'hFEC3;
    16'd46580: out <= 16'hFF17;    16'd46581: out <= 16'hFEDA;    16'd46582: out <= 16'hFF45;    16'd46583: out <= 16'h009F;
    16'd46584: out <= 16'h0963;    16'd46585: out <= 16'h038F;    16'd46586: out <= 16'h0171;    16'd46587: out <= 16'hFEB6;
    16'd46588: out <= 16'hFC84;    16'd46589: out <= 16'hFA46;    16'd46590: out <= 16'h0213;    16'd46591: out <= 16'hFF81;
    16'd46592: out <= 16'hFEAE;    16'd46593: out <= 16'hFD8D;    16'd46594: out <= 16'h02BF;    16'd46595: out <= 16'hFD19;
    16'd46596: out <= 16'h02B9;    16'd46597: out <= 16'hF9FA;    16'd46598: out <= 16'h0126;    16'd46599: out <= 16'h03DF;
    16'd46600: out <= 16'hF873;    16'd46601: out <= 16'hFE7D;    16'd46602: out <= 16'hFC67;    16'd46603: out <= 16'h0204;
    16'd46604: out <= 16'hFB81;    16'd46605: out <= 16'h06FC;    16'd46606: out <= 16'h02BF;    16'd46607: out <= 16'h0458;
    16'd46608: out <= 16'hF893;    16'd46609: out <= 16'h00E4;    16'd46610: out <= 16'h0092;    16'd46611: out <= 16'h0283;
    16'd46612: out <= 16'h034F;    16'd46613: out <= 16'h0281;    16'd46614: out <= 16'h00D0;    16'd46615: out <= 16'hFC40;
    16'd46616: out <= 16'h0005;    16'd46617: out <= 16'h0148;    16'd46618: out <= 16'h01F1;    16'd46619: out <= 16'hFFED;
    16'd46620: out <= 16'hFBA5;    16'd46621: out <= 16'hFD10;    16'd46622: out <= 16'hFE02;    16'd46623: out <= 16'h030B;
    16'd46624: out <= 16'hFF4B;    16'd46625: out <= 16'h000B;    16'd46626: out <= 16'h0362;    16'd46627: out <= 16'hFCCD;
    16'd46628: out <= 16'h00EE;    16'd46629: out <= 16'hFFBD;    16'd46630: out <= 16'h0714;    16'd46631: out <= 16'hFF97;
    16'd46632: out <= 16'h011B;    16'd46633: out <= 16'h04FA;    16'd46634: out <= 16'h0201;    16'd46635: out <= 16'h0345;
    16'd46636: out <= 16'h049B;    16'd46637: out <= 16'h04D9;    16'd46638: out <= 16'h0E8D;    16'd46639: out <= 16'h0CA8;
    16'd46640: out <= 16'h062B;    16'd46641: out <= 16'hFFEA;    16'd46642: out <= 16'h07C6;    16'd46643: out <= 16'h00B5;
    16'd46644: out <= 16'hFAB6;    16'd46645: out <= 16'h04DE;    16'd46646: out <= 16'h014B;    16'd46647: out <= 16'h0891;
    16'd46648: out <= 16'h02E0;    16'd46649: out <= 16'h0308;    16'd46650: out <= 16'h08EA;    16'd46651: out <= 16'hFFE0;
    16'd46652: out <= 16'h06FB;    16'd46653: out <= 16'h0427;    16'd46654: out <= 16'hFFBD;    16'd46655: out <= 16'h0347;
    16'd46656: out <= 16'h0982;    16'd46657: out <= 16'h095D;    16'd46658: out <= 16'h031B;    16'd46659: out <= 16'h0160;
    16'd46660: out <= 16'h0080;    16'd46661: out <= 16'h019A;    16'd46662: out <= 16'hFC02;    16'd46663: out <= 16'hFF3A;
    16'd46664: out <= 16'hFE3A;    16'd46665: out <= 16'h02C1;    16'd46666: out <= 16'hFDBF;    16'd46667: out <= 16'h0001;
    16'd46668: out <= 16'hFF62;    16'd46669: out <= 16'h02A4;    16'd46670: out <= 16'hFF49;    16'd46671: out <= 16'h000D;
    16'd46672: out <= 16'hFE7C;    16'd46673: out <= 16'h04B8;    16'd46674: out <= 16'hFF3B;    16'd46675: out <= 16'h001F;
    16'd46676: out <= 16'h048D;    16'd46677: out <= 16'hFFC0;    16'd46678: out <= 16'h00C5;    16'd46679: out <= 16'h00E9;
    16'd46680: out <= 16'hFD19;    16'd46681: out <= 16'hFC8A;    16'd46682: out <= 16'hFEF3;    16'd46683: out <= 16'hFA2D;
    16'd46684: out <= 16'h032D;    16'd46685: out <= 16'h0466;    16'd46686: out <= 16'hFD29;    16'd46687: out <= 16'h00E0;
    16'd46688: out <= 16'hFD70;    16'd46689: out <= 16'h0549;    16'd46690: out <= 16'hFF61;    16'd46691: out <= 16'hFE7A;
    16'd46692: out <= 16'hFF15;    16'd46693: out <= 16'h03F8;    16'd46694: out <= 16'hFE6C;    16'd46695: out <= 16'hFC18;
    16'd46696: out <= 16'hF95A;    16'd46697: out <= 16'hFFCC;    16'd46698: out <= 16'hFD8F;    16'd46699: out <= 16'hFF8D;
    16'd46700: out <= 16'hFE86;    16'd46701: out <= 16'h0055;    16'd46702: out <= 16'hFC63;    16'd46703: out <= 16'h0095;
    16'd46704: out <= 16'hF95E;    16'd46705: out <= 16'hFF47;    16'd46706: out <= 16'hFD88;    16'd46707: out <= 16'h037E;
    16'd46708: out <= 16'h01C0;    16'd46709: out <= 16'h0069;    16'd46710: out <= 16'h0736;    16'd46711: out <= 16'hFC8D;
    16'd46712: out <= 16'h00AF;    16'd46713: out <= 16'h01DD;    16'd46714: out <= 16'h0135;    16'd46715: out <= 16'h01CE;
    16'd46716: out <= 16'hFEE2;    16'd46717: out <= 16'h0208;    16'd46718: out <= 16'hFB80;    16'd46719: out <= 16'hF773;
    16'd46720: out <= 16'hFFD1;    16'd46721: out <= 16'hF89A;    16'd46722: out <= 16'hFDC9;    16'd46723: out <= 16'h03C6;
    16'd46724: out <= 16'hFD1A;    16'd46725: out <= 16'hF6CB;    16'd46726: out <= 16'hFEB4;    16'd46727: out <= 16'h0213;
    16'd46728: out <= 16'hFDF0;    16'd46729: out <= 16'h0739;    16'd46730: out <= 16'h05C5;    16'd46731: out <= 16'hFEF3;
    16'd46732: out <= 16'h0592;    16'd46733: out <= 16'h03B1;    16'd46734: out <= 16'h0726;    16'd46735: out <= 16'hFDE2;
    16'd46736: out <= 16'h0080;    16'd46737: out <= 16'h0091;    16'd46738: out <= 16'h05DE;    16'd46739: out <= 16'h068B;
    16'd46740: out <= 16'h0980;    16'd46741: out <= 16'h06E0;    16'd46742: out <= 16'h018B;    16'd46743: out <= 16'h0571;
    16'd46744: out <= 16'h07E4;    16'd46745: out <= 16'h0869;    16'd46746: out <= 16'h029A;    16'd46747: out <= 16'hFF13;
    16'd46748: out <= 16'h05D5;    16'd46749: out <= 16'hFDB6;    16'd46750: out <= 16'h048B;    16'd46751: out <= 16'h09B0;
    16'd46752: out <= 16'h038C;    16'd46753: out <= 16'hFD67;    16'd46754: out <= 16'h050A;    16'd46755: out <= 16'h025E;
    16'd46756: out <= 16'h0546;    16'd46757: out <= 16'h0056;    16'd46758: out <= 16'h0241;    16'd46759: out <= 16'h0749;
    16'd46760: out <= 16'h01F9;    16'd46761: out <= 16'h077D;    16'd46762: out <= 16'h02BE;    16'd46763: out <= 16'h0A1C;
    16'd46764: out <= 16'h04A6;    16'd46765: out <= 16'h0353;    16'd46766: out <= 16'h06A2;    16'd46767: out <= 16'h00BC;
    16'd46768: out <= 16'h043D;    16'd46769: out <= 16'h052B;    16'd46770: out <= 16'h0885;    16'd46771: out <= 16'h02BC;
    16'd46772: out <= 16'hFFD2;    16'd46773: out <= 16'hFEEF;    16'd46774: out <= 16'h0509;    16'd46775: out <= 16'h076F;
    16'd46776: out <= 16'h07C1;    16'd46777: out <= 16'h00C1;    16'd46778: out <= 16'h0FAA;    16'd46779: out <= 16'h05D2;
    16'd46780: out <= 16'h043E;    16'd46781: out <= 16'h0728;    16'd46782: out <= 16'h087D;    16'd46783: out <= 16'h058A;
    16'd46784: out <= 16'h069A;    16'd46785: out <= 16'h07D3;    16'd46786: out <= 16'h03D5;    16'd46787: out <= 16'h04AE;
    16'd46788: out <= 16'h0070;    16'd46789: out <= 16'hFDF1;    16'd46790: out <= 16'h00E4;    16'd46791: out <= 16'hFD79;
    16'd46792: out <= 16'h01D7;    16'd46793: out <= 16'h0101;    16'd46794: out <= 16'h02C2;    16'd46795: out <= 16'h02A8;
    16'd46796: out <= 16'h01EB;    16'd46797: out <= 16'hFAE3;    16'd46798: out <= 16'hFFF5;    16'd46799: out <= 16'hFC8B;
    16'd46800: out <= 16'hFD6A;    16'd46801: out <= 16'hFD49;    16'd46802: out <= 16'h06EA;    16'd46803: out <= 16'hFEF9;
    16'd46804: out <= 16'h0195;    16'd46805: out <= 16'hF985;    16'd46806: out <= 16'hF92B;    16'd46807: out <= 16'h02FD;
    16'd46808: out <= 16'hF9D4;    16'd46809: out <= 16'hFF6F;    16'd46810: out <= 16'h0348;    16'd46811: out <= 16'hFE82;
    16'd46812: out <= 16'hFC19;    16'd46813: out <= 16'hFFB4;    16'd46814: out <= 16'hFEBD;    16'd46815: out <= 16'hFDD1;
    16'd46816: out <= 16'hFC35;    16'd46817: out <= 16'h04EC;    16'd46818: out <= 16'h016D;    16'd46819: out <= 16'h072D;
    16'd46820: out <= 16'hFE19;    16'd46821: out <= 16'h0465;    16'd46822: out <= 16'hF811;    16'd46823: out <= 16'h009D;
    16'd46824: out <= 16'h019A;    16'd46825: out <= 16'hF6C9;    16'd46826: out <= 16'h02EA;    16'd46827: out <= 16'hFD85;
    16'd46828: out <= 16'h0597;    16'd46829: out <= 16'h0938;    16'd46830: out <= 16'h0304;    16'd46831: out <= 16'h01E8;
    16'd46832: out <= 16'h020F;    16'd46833: out <= 16'hFDE6;    16'd46834: out <= 16'h026F;    16'd46835: out <= 16'hFB8B;
    16'd46836: out <= 16'h00E7;    16'd46837: out <= 16'hFD88;    16'd46838: out <= 16'h04C1;    16'd46839: out <= 16'h0274;
    16'd46840: out <= 16'hFE4E;    16'd46841: out <= 16'h002B;    16'd46842: out <= 16'h032A;    16'd46843: out <= 16'hFDB5;
    16'd46844: out <= 16'hF9DE;    16'd46845: out <= 16'hFBDF;    16'd46846: out <= 16'h033B;    16'd46847: out <= 16'h00D7;
    16'd46848: out <= 16'hFE00;    16'd46849: out <= 16'hFA40;    16'd46850: out <= 16'h00BA;    16'd46851: out <= 16'h00BA;
    16'd46852: out <= 16'hFE2B;    16'd46853: out <= 16'h069B;    16'd46854: out <= 16'hFC0D;    16'd46855: out <= 16'hFC5E;
    16'd46856: out <= 16'h011A;    16'd46857: out <= 16'h07AB;    16'd46858: out <= 16'h020B;    16'd46859: out <= 16'h069D;
    16'd46860: out <= 16'hFF1C;    16'd46861: out <= 16'h0557;    16'd46862: out <= 16'hFD4F;    16'd46863: out <= 16'hFB57;
    16'd46864: out <= 16'h0407;    16'd46865: out <= 16'hFF99;    16'd46866: out <= 16'hFFC1;    16'd46867: out <= 16'h00CC;
    16'd46868: out <= 16'h03ED;    16'd46869: out <= 16'hFFD2;    16'd46870: out <= 16'h07E2;    16'd46871: out <= 16'hF8E5;
    16'd46872: out <= 16'h01C8;    16'd46873: out <= 16'hFDFD;    16'd46874: out <= 16'h042A;    16'd46875: out <= 16'hFF03;
    16'd46876: out <= 16'h0369;    16'd46877: out <= 16'hF9D7;    16'd46878: out <= 16'h0439;    16'd46879: out <= 16'hFF94;
    16'd46880: out <= 16'h0103;    16'd46881: out <= 16'h0462;    16'd46882: out <= 16'hFD5B;    16'd46883: out <= 16'h004A;
    16'd46884: out <= 16'hF9C8;    16'd46885: out <= 16'h032B;    16'd46886: out <= 16'h05E9;    16'd46887: out <= 16'h06AC;
    16'd46888: out <= 16'h0CFB;    16'd46889: out <= 16'hFF84;    16'd46890: out <= 16'h0C30;    16'd46891: out <= 16'hFFA7;
    16'd46892: out <= 16'h036B;    16'd46893: out <= 16'h052A;    16'd46894: out <= 16'h0A2C;    16'd46895: out <= 16'h00F3;
    16'd46896: out <= 16'h0771;    16'd46897: out <= 16'h0520;    16'd46898: out <= 16'h08EF;    16'd46899: out <= 16'h0045;
    16'd46900: out <= 16'h0769;    16'd46901: out <= 16'h02E4;    16'd46902: out <= 16'h08DF;    16'd46903: out <= 16'h0B07;
    16'd46904: out <= 16'h05F7;    16'd46905: out <= 16'h0483;    16'd46906: out <= 16'h066F;    16'd46907: out <= 16'h075D;
    16'd46908: out <= 16'h02D4;    16'd46909: out <= 16'h0226;    16'd46910: out <= 16'hFE48;    16'd46911: out <= 16'h056A;
    16'd46912: out <= 16'h0693;    16'd46913: out <= 16'hFF10;    16'd46914: out <= 16'hFEBF;    16'd46915: out <= 16'h0178;
    16'd46916: out <= 16'h09CB;    16'd46917: out <= 16'h0387;    16'd46918: out <= 16'h006B;    16'd46919: out <= 16'h069E;
    16'd46920: out <= 16'hFF20;    16'd46921: out <= 16'h060A;    16'd46922: out <= 16'hFD8F;    16'd46923: out <= 16'hFCE7;
    16'd46924: out <= 16'hF7C5;    16'd46925: out <= 16'hFCD7;    16'd46926: out <= 16'hFE1A;    16'd46927: out <= 16'h024F;
    16'd46928: out <= 16'hFABD;    16'd46929: out <= 16'hFE79;    16'd46930: out <= 16'h002A;    16'd46931: out <= 16'hFF6D;
    16'd46932: out <= 16'hFDE8;    16'd46933: out <= 16'h03DB;    16'd46934: out <= 16'h02A3;    16'd46935: out <= 16'hFE5F;
    16'd46936: out <= 16'h02E0;    16'd46937: out <= 16'h0645;    16'd46938: out <= 16'hFD31;    16'd46939: out <= 16'hFD7D;
    16'd46940: out <= 16'h048E;    16'd46941: out <= 16'h0496;    16'd46942: out <= 16'hFBF8;    16'd46943: out <= 16'h0107;
    16'd46944: out <= 16'h0084;    16'd46945: out <= 16'hFF22;    16'd46946: out <= 16'hF9E5;    16'd46947: out <= 16'hF9B1;
    16'd46948: out <= 16'h07C0;    16'd46949: out <= 16'hFF8C;    16'd46950: out <= 16'hFED8;    16'd46951: out <= 16'hFA2A;
    16'd46952: out <= 16'h0434;    16'd46953: out <= 16'h02FD;    16'd46954: out <= 16'h0550;    16'd46955: out <= 16'hFF59;
    16'd46956: out <= 16'hFB1D;    16'd46957: out <= 16'h049A;    16'd46958: out <= 16'hFDE2;    16'd46959: out <= 16'h062E;
    16'd46960: out <= 16'hFDBA;    16'd46961: out <= 16'h011E;    16'd46962: out <= 16'h009E;    16'd46963: out <= 16'h005C;
    16'd46964: out <= 16'h00C6;    16'd46965: out <= 16'hFCFC;    16'd46966: out <= 16'h026D;    16'd46967: out <= 16'h023E;
    16'd46968: out <= 16'hFEBB;    16'd46969: out <= 16'hFF81;    16'd46970: out <= 16'hFEEA;    16'd46971: out <= 16'hFF6C;
    16'd46972: out <= 16'hFCD8;    16'd46973: out <= 16'hFDA2;    16'd46974: out <= 16'h040D;    16'd46975: out <= 16'h01A3;
    16'd46976: out <= 16'h010A;    16'd46977: out <= 16'hFF4F;    16'd46978: out <= 16'h024B;    16'd46979: out <= 16'hFC59;
    16'd46980: out <= 16'h03DD;    16'd46981: out <= 16'hFD03;    16'd46982: out <= 16'h0459;    16'd46983: out <= 16'h01D0;
    16'd46984: out <= 16'h01B1;    16'd46985: out <= 16'hFE6D;    16'd46986: out <= 16'h0106;    16'd46987: out <= 16'hF9E7;
    16'd46988: out <= 16'h0714;    16'd46989: out <= 16'h08E0;    16'd46990: out <= 16'h0104;    16'd46991: out <= 16'hFE60;
    16'd46992: out <= 16'h0875;    16'd46993: out <= 16'h02F7;    16'd46994: out <= 16'h0509;    16'd46995: out <= 16'h01F2;
    16'd46996: out <= 16'h03AF;    16'd46997: out <= 16'h08E1;    16'd46998: out <= 16'h0554;    16'd46999: out <= 16'h0764;
    16'd47000: out <= 16'h0432;    16'd47001: out <= 16'h01D9;    16'd47002: out <= 16'h0561;    16'd47003: out <= 16'h04A7;
    16'd47004: out <= 16'h06CF;    16'd47005: out <= 16'hFF24;    16'd47006: out <= 16'h007E;    16'd47007: out <= 16'h0719;
    16'd47008: out <= 16'h058A;    16'd47009: out <= 16'h0060;    16'd47010: out <= 16'h04D0;    16'd47011: out <= 16'h0557;
    16'd47012: out <= 16'hFF23;    16'd47013: out <= 16'h0617;    16'd47014: out <= 16'h04C7;    16'd47015: out <= 16'h0ED0;
    16'd47016: out <= 16'h01F7;    16'd47017: out <= 16'hFEF4;    16'd47018: out <= 16'hFF0F;    16'd47019: out <= 16'h02CF;
    16'd47020: out <= 16'h00E3;    16'd47021: out <= 16'h0502;    16'd47022: out <= 16'h0708;    16'd47023: out <= 16'h02FF;
    16'd47024: out <= 16'h00BC;    16'd47025: out <= 16'h02A2;    16'd47026: out <= 16'h0456;    16'd47027: out <= 16'hFABD;
    16'd47028: out <= 16'h03DE;    16'd47029: out <= 16'h072F;    16'd47030: out <= 16'h0526;    16'd47031: out <= 16'h0900;
    16'd47032: out <= 16'hFC1C;    16'd47033: out <= 16'h0450;    16'd47034: out <= 16'h050D;    16'd47035: out <= 16'h0573;
    16'd47036: out <= 16'h0200;    16'd47037: out <= 16'h005E;    16'd47038: out <= 16'h0885;    16'd47039: out <= 16'h0166;
    16'd47040: out <= 16'h007E;    16'd47041: out <= 16'h0270;    16'd47042: out <= 16'h08D2;    16'd47043: out <= 16'h0564;
    16'd47044: out <= 16'hFEF7;    16'd47045: out <= 16'h0528;    16'd47046: out <= 16'h00EE;    16'd47047: out <= 16'h048B;
    16'd47048: out <= 16'h04C3;    16'd47049: out <= 16'h012A;    16'd47050: out <= 16'h01AE;    16'd47051: out <= 16'hFFF2;
    16'd47052: out <= 16'hFDB6;    16'd47053: out <= 16'hFF04;    16'd47054: out <= 16'hFA92;    16'd47055: out <= 16'hFCE6;
    16'd47056: out <= 16'hFC8D;    16'd47057: out <= 16'h0406;    16'd47058: out <= 16'hFEBF;    16'd47059: out <= 16'h02D8;
    16'd47060: out <= 16'hFE07;    16'd47061: out <= 16'h032C;    16'd47062: out <= 16'h02AD;    16'd47063: out <= 16'hFDF7;
    16'd47064: out <= 16'hFC9D;    16'd47065: out <= 16'hFC84;    16'd47066: out <= 16'h0007;    16'd47067: out <= 16'hFEF8;
    16'd47068: out <= 16'h006B;    16'd47069: out <= 16'h0500;    16'd47070: out <= 16'h0945;    16'd47071: out <= 16'h045D;
    16'd47072: out <= 16'hFD85;    16'd47073: out <= 16'h0020;    16'd47074: out <= 16'hF73D;    16'd47075: out <= 16'h0457;
    16'd47076: out <= 16'h011A;    16'd47077: out <= 16'h00DC;    16'd47078: out <= 16'hFEF9;    16'd47079: out <= 16'hFF77;
    16'd47080: out <= 16'hF5F8;    16'd47081: out <= 16'h0195;    16'd47082: out <= 16'hFF6C;    16'd47083: out <= 16'h0162;
    16'd47084: out <= 16'h02A2;    16'd47085: out <= 16'h075F;    16'd47086: out <= 16'hFF89;    16'd47087: out <= 16'hFDBE;
    16'd47088: out <= 16'h00B9;    16'd47089: out <= 16'hF956;    16'd47090: out <= 16'hF93F;    16'd47091: out <= 16'h0245;
    16'd47092: out <= 16'hF718;    16'd47093: out <= 16'h00E6;    16'd47094: out <= 16'hF95B;    16'd47095: out <= 16'hFD9E;
    16'd47096: out <= 16'hFC0A;    16'd47097: out <= 16'h0129;    16'd47098: out <= 16'hFFC7;    16'd47099: out <= 16'h0123;
    16'd47100: out <= 16'h07B1;    16'd47101: out <= 16'hFE9C;    16'd47102: out <= 16'hF8E8;    16'd47103: out <= 16'h01A0;
    16'd47104: out <= 16'hF7B0;    16'd47105: out <= 16'hFDD2;    16'd47106: out <= 16'hFEF0;    16'd47107: out <= 16'h0363;
    16'd47108: out <= 16'h021F;    16'd47109: out <= 16'h0442;    16'd47110: out <= 16'h0284;    16'd47111: out <= 16'h026F;
    16'd47112: out <= 16'hFFFB;    16'd47113: out <= 16'h0121;    16'd47114: out <= 16'hF974;    16'd47115: out <= 16'h04B6;
    16'd47116: out <= 16'h00EE;    16'd47117: out <= 16'hFA76;    16'd47118: out <= 16'hF925;    16'd47119: out <= 16'h00FE;
    16'd47120: out <= 16'hFE31;    16'd47121: out <= 16'h00F6;    16'd47122: out <= 16'h03E4;    16'd47123: out <= 16'h0842;
    16'd47124: out <= 16'h07AD;    16'd47125: out <= 16'hFE8C;    16'd47126: out <= 16'hFD74;    16'd47127: out <= 16'h0776;
    16'd47128: out <= 16'h02A5;    16'd47129: out <= 16'h00BC;    16'd47130: out <= 16'h0343;    16'd47131: out <= 16'h0033;
    16'd47132: out <= 16'hFD46;    16'd47133: out <= 16'hFC63;    16'd47134: out <= 16'hFDF3;    16'd47135: out <= 16'hFDD2;
    16'd47136: out <= 16'h0277;    16'd47137: out <= 16'h035E;    16'd47138: out <= 16'h01F2;    16'd47139: out <= 16'hFC0C;
    16'd47140: out <= 16'h0114;    16'd47141: out <= 16'h070C;    16'd47142: out <= 16'hFF2A;    16'd47143: out <= 16'h0644;
    16'd47144: out <= 16'h075C;    16'd47145: out <= 16'h0F10;    16'd47146: out <= 16'h06DE;    16'd47147: out <= 16'hFE9D;
    16'd47148: out <= 16'h0ADF;    16'd47149: out <= 16'h0269;    16'd47150: out <= 16'h04C5;    16'd47151: out <= 16'h05C4;
    16'd47152: out <= 16'h0001;    16'd47153: out <= 16'h0531;    16'd47154: out <= 16'h0148;    16'd47155: out <= 16'h0655;
    16'd47156: out <= 16'h0636;    16'd47157: out <= 16'h01B2;    16'd47158: out <= 16'h107B;    16'd47159: out <= 16'hFD17;
    16'd47160: out <= 16'h035F;    16'd47161: out <= 16'hFE75;    16'd47162: out <= 16'h082C;    16'd47163: out <= 16'h0548;
    16'd47164: out <= 16'h0876;    16'd47165: out <= 16'h05C4;    16'd47166: out <= 16'hFE98;    16'd47167: out <= 16'h018E;
    16'd47168: out <= 16'h045A;    16'd47169: out <= 16'h0148;    16'd47170: out <= 16'h0967;    16'd47171: out <= 16'h094A;
    16'd47172: out <= 16'h03A2;    16'd47173: out <= 16'hFDFF;    16'd47174: out <= 16'h054E;    16'd47175: out <= 16'h0326;
    16'd47176: out <= 16'h00CC;    16'd47177: out <= 16'h02A0;    16'd47178: out <= 16'h0144;    16'd47179: out <= 16'h01C4;
    16'd47180: out <= 16'h015E;    16'd47181: out <= 16'hFFBD;    16'd47182: out <= 16'h005D;    16'd47183: out <= 16'h027C;
    16'd47184: out <= 16'h002E;    16'd47185: out <= 16'hFEE1;    16'd47186: out <= 16'hFDDD;    16'd47187: out <= 16'h057F;
    16'd47188: out <= 16'h01A7;    16'd47189: out <= 16'h0198;    16'd47190: out <= 16'hFE5D;    16'd47191: out <= 16'hFA77;
    16'd47192: out <= 16'h0380;    16'd47193: out <= 16'hFF7E;    16'd47194: out <= 16'h05EE;    16'd47195: out <= 16'h0235;
    16'd47196: out <= 16'h0541;    16'd47197: out <= 16'h022F;    16'd47198: out <= 16'h0768;    16'd47199: out <= 16'h0A1F;
    16'd47200: out <= 16'h0399;    16'd47201: out <= 16'hFCEB;    16'd47202: out <= 16'h0595;    16'd47203: out <= 16'h04A8;
    16'd47204: out <= 16'hFCE5;    16'd47205: out <= 16'h0668;    16'd47206: out <= 16'h020A;    16'd47207: out <= 16'h004A;
    16'd47208: out <= 16'hFDF4;    16'd47209: out <= 16'hFB99;    16'd47210: out <= 16'hFD75;    16'd47211: out <= 16'h0036;
    16'd47212: out <= 16'hFA1B;    16'd47213: out <= 16'h06FF;    16'd47214: out <= 16'hFEBF;    16'd47215: out <= 16'hFA33;
    16'd47216: out <= 16'hFEDC;    16'd47217: out <= 16'hFF04;    16'd47218: out <= 16'hFF2B;    16'd47219: out <= 16'hFFF1;
    16'd47220: out <= 16'hFC68;    16'd47221: out <= 16'h01EC;    16'd47222: out <= 16'hFEA6;    16'd47223: out <= 16'hFE0D;
    16'd47224: out <= 16'h06F3;    16'd47225: out <= 16'h0031;    16'd47226: out <= 16'hFBB8;    16'd47227: out <= 16'hFEF5;
    16'd47228: out <= 16'hFDF0;    16'd47229: out <= 16'hF6B6;    16'd47230: out <= 16'hFA7C;    16'd47231: out <= 16'h065A;
    16'd47232: out <= 16'hF98C;    16'd47233: out <= 16'hFF92;    16'd47234: out <= 16'hFEB7;    16'd47235: out <= 16'hFD24;
    16'd47236: out <= 16'h0101;    16'd47237: out <= 16'h01E1;    16'd47238: out <= 16'hFBFC;    16'd47239: out <= 16'h0248;
    16'd47240: out <= 16'hFC02;    16'd47241: out <= 16'h0051;    16'd47242: out <= 16'h00E7;    16'd47243: out <= 16'hFF35;
    16'd47244: out <= 16'hFF5C;    16'd47245: out <= 16'hFA9D;    16'd47246: out <= 16'hFF14;    16'd47247: out <= 16'hFF97;
    16'd47248: out <= 16'h0933;    16'd47249: out <= 16'hFFD1;    16'd47250: out <= 16'h0492;    16'd47251: out <= 16'h0392;
    16'd47252: out <= 16'h094D;    16'd47253: out <= 16'h024A;    16'd47254: out <= 16'h002D;    16'd47255: out <= 16'h02F4;
    16'd47256: out <= 16'h003B;    16'd47257: out <= 16'h031B;    16'd47258: out <= 16'h057D;    16'd47259: out <= 16'hFEE7;
    16'd47260: out <= 16'h0452;    16'd47261: out <= 16'h040F;    16'd47262: out <= 16'h0004;    16'd47263: out <= 16'h0580;
    16'd47264: out <= 16'h0557;    16'd47265: out <= 16'h083B;    16'd47266: out <= 16'hFFB1;    16'd47267: out <= 16'h0357;
    16'd47268: out <= 16'h0403;    16'd47269: out <= 16'h003F;    16'd47270: out <= 16'h0607;    16'd47271: out <= 16'h01BC;
    16'd47272: out <= 16'hFF59;    16'd47273: out <= 16'hFEAB;    16'd47274: out <= 16'h05D7;    16'd47275: out <= 16'h0430;
    16'd47276: out <= 16'hFB68;    16'd47277: out <= 16'h0699;    16'd47278: out <= 16'hFE11;    16'd47279: out <= 16'h08C6;
    16'd47280: out <= 16'h0350;    16'd47281: out <= 16'hFEE4;    16'd47282: out <= 16'h04A0;    16'd47283: out <= 16'h01D0;
    16'd47284: out <= 16'h0219;    16'd47285: out <= 16'h0744;    16'd47286: out <= 16'hFF2F;    16'd47287: out <= 16'h0094;
    16'd47288: out <= 16'h06A2;    16'd47289: out <= 16'h0581;    16'd47290: out <= 16'h086A;    16'd47291: out <= 16'h055D;
    16'd47292: out <= 16'h00B3;    16'd47293: out <= 16'h0483;    16'd47294: out <= 16'h0339;    16'd47295: out <= 16'h0641;
    16'd47296: out <= 16'h07A7;    16'd47297: out <= 16'h00FB;    16'd47298: out <= 16'h0917;    16'd47299: out <= 16'h0072;
    16'd47300: out <= 16'h0181;    16'd47301: out <= 16'h0B1C;    16'd47302: out <= 16'h090D;    16'd47303: out <= 16'h01B9;
    16'd47304: out <= 16'hFF70;    16'd47305: out <= 16'hFF17;    16'd47306: out <= 16'hFC3E;    16'd47307: out <= 16'hFD34;
    16'd47308: out <= 16'hFCCF;    16'd47309: out <= 16'h04A8;    16'd47310: out <= 16'h066D;    16'd47311: out <= 16'h049D;
    16'd47312: out <= 16'hFB30;    16'd47313: out <= 16'h042E;    16'd47314: out <= 16'hFEB7;    16'd47315: out <= 16'h04B3;
    16'd47316: out <= 16'hFAA5;    16'd47317: out <= 16'h090F;    16'd47318: out <= 16'h00FF;    16'd47319: out <= 16'hFE33;
    16'd47320: out <= 16'h02EB;    16'd47321: out <= 16'hFDC0;    16'd47322: out <= 16'hFD3F;    16'd47323: out <= 16'hFFF8;
    16'd47324: out <= 16'hFDDC;    16'd47325: out <= 16'h0527;    16'd47326: out <= 16'hFC44;    16'd47327: out <= 16'h066C;
    16'd47328: out <= 16'h044F;    16'd47329: out <= 16'h0616;    16'd47330: out <= 16'hFF8E;    16'd47331: out <= 16'hFE5E;
    16'd47332: out <= 16'hFE90;    16'd47333: out <= 16'h00A0;    16'd47334: out <= 16'h080E;    16'd47335: out <= 16'h01BB;
    16'd47336: out <= 16'hFD24;    16'd47337: out <= 16'h002F;    16'd47338: out <= 16'h0397;    16'd47339: out <= 16'hFCB3;
    16'd47340: out <= 16'hF9C0;    16'd47341: out <= 16'hFFF2;    16'd47342: out <= 16'h01C9;    16'd47343: out <= 16'h0807;
    16'd47344: out <= 16'hFEFB;    16'd47345: out <= 16'h0025;    16'd47346: out <= 16'h003E;    16'd47347: out <= 16'hFD7F;
    16'd47348: out <= 16'h0079;    16'd47349: out <= 16'hFFA9;    16'd47350: out <= 16'h05F6;    16'd47351: out <= 16'h00AE;
    16'd47352: out <= 16'hFD4C;    16'd47353: out <= 16'hFFB5;    16'd47354: out <= 16'h02D7;    16'd47355: out <= 16'hFD07;
    16'd47356: out <= 16'h01A5;    16'd47357: out <= 16'h04CD;    16'd47358: out <= 16'h0269;    16'd47359: out <= 16'h0092;
    16'd47360: out <= 16'h01CA;    16'd47361: out <= 16'h0167;    16'd47362: out <= 16'h038E;    16'd47363: out <= 16'hFB6E;
    16'd47364: out <= 16'h091D;    16'd47365: out <= 16'h02D4;    16'd47366: out <= 16'h017C;    16'd47367: out <= 16'hFEA4;
    16'd47368: out <= 16'hFF82;    16'd47369: out <= 16'hFFB5;    16'd47370: out <= 16'hFD2D;    16'd47371: out <= 16'hFB1D;
    16'd47372: out <= 16'h0319;    16'd47373: out <= 16'h02CD;    16'd47374: out <= 16'hF8DA;    16'd47375: out <= 16'hFAD4;
    16'd47376: out <= 16'h033C;    16'd47377: out <= 16'hFE18;    16'd47378: out <= 16'h026D;    16'd47379: out <= 16'h00C3;
    16'd47380: out <= 16'h089D;    16'd47381: out <= 16'hFBFB;    16'd47382: out <= 16'hF881;    16'd47383: out <= 16'h0167;
    16'd47384: out <= 16'hFFBC;    16'd47385: out <= 16'hFDB5;    16'd47386: out <= 16'hFBDE;    16'd47387: out <= 16'h028D;
    16'd47388: out <= 16'hFEE7;    16'd47389: out <= 16'h033C;    16'd47390: out <= 16'hFFFD;    16'd47391: out <= 16'h0600;
    16'd47392: out <= 16'h072C;    16'd47393: out <= 16'hFEA6;    16'd47394: out <= 16'h05BA;    16'd47395: out <= 16'h0443;
    16'd47396: out <= 16'hFE23;    16'd47397: out <= 16'hFE7F;    16'd47398: out <= 16'h021F;    16'd47399: out <= 16'h05C5;
    16'd47400: out <= 16'hFD3B;    16'd47401: out <= 16'h03D3;    16'd47402: out <= 16'h0625;    16'd47403: out <= 16'h044F;
    16'd47404: out <= 16'h01D6;    16'd47405: out <= 16'h03B6;    16'd47406: out <= 16'h0688;    16'd47407: out <= 16'hFE53;
    16'd47408: out <= 16'h0397;    16'd47409: out <= 16'h049A;    16'd47410: out <= 16'hFFF5;    16'd47411: out <= 16'h060E;
    16'd47412: out <= 16'hFEA3;    16'd47413: out <= 16'h094A;    16'd47414: out <= 16'h0588;    16'd47415: out <= 16'hFE13;
    16'd47416: out <= 16'h0291;    16'd47417: out <= 16'h024B;    16'd47418: out <= 16'h03D3;    16'd47419: out <= 16'h0476;
    16'd47420: out <= 16'h07A0;    16'd47421: out <= 16'h0510;    16'd47422: out <= 16'h03BE;    16'd47423: out <= 16'h0116;
    16'd47424: out <= 16'hFC97;    16'd47425: out <= 16'h01C8;    16'd47426: out <= 16'h0760;    16'd47427: out <= 16'h0575;
    16'd47428: out <= 16'h084B;    16'd47429: out <= 16'h0738;    16'd47430: out <= 16'h0237;    16'd47431: out <= 16'hFEA4;
    16'd47432: out <= 16'h003E;    16'd47433: out <= 16'hFF7A;    16'd47434: out <= 16'hFAD4;    16'd47435: out <= 16'hFC9E;
    16'd47436: out <= 16'h001B;    16'd47437: out <= 16'h01E1;    16'd47438: out <= 16'hFABD;    16'd47439: out <= 16'hFAB6;
    16'd47440: out <= 16'hFAFB;    16'd47441: out <= 16'h0D6F;    16'd47442: out <= 16'h041E;    16'd47443: out <= 16'h0096;
    16'd47444: out <= 16'h0353;    16'd47445: out <= 16'h0503;    16'd47446: out <= 16'h0203;    16'd47447: out <= 16'h008E;
    16'd47448: out <= 16'h0201;    16'd47449: out <= 16'h07D1;    16'd47450: out <= 16'h0615;    16'd47451: out <= 16'h01E6;
    16'd47452: out <= 16'h02A8;    16'd47453: out <= 16'h073D;    16'd47454: out <= 16'h043E;    16'd47455: out <= 16'hFE1A;
    16'd47456: out <= 16'h02E6;    16'd47457: out <= 16'hFDF2;    16'd47458: out <= 16'h00D4;    16'd47459: out <= 16'h027F;
    16'd47460: out <= 16'hFEA1;    16'd47461: out <= 16'hFE90;    16'd47462: out <= 16'hF9BC;    16'd47463: out <= 16'h02F4;
    16'd47464: out <= 16'hFE76;    16'd47465: out <= 16'hFD86;    16'd47466: out <= 16'h02E1;    16'd47467: out <= 16'h01B2;
    16'd47468: out <= 16'hF8CE;    16'd47469: out <= 16'hF530;    16'd47470: out <= 16'hF37C;    16'd47471: out <= 16'hFF8F;
    16'd47472: out <= 16'hFC49;    16'd47473: out <= 16'h0553;    16'd47474: out <= 16'hFCD1;    16'd47475: out <= 16'hFC66;
    16'd47476: out <= 16'hFED8;    16'd47477: out <= 16'hFB77;    16'd47478: out <= 16'h0006;    16'd47479: out <= 16'hFF40;
    16'd47480: out <= 16'h0993;    16'd47481: out <= 16'hFAAB;    16'd47482: out <= 16'hFD7F;    16'd47483: out <= 16'h01FA;
    16'd47484: out <= 16'h0231;    16'd47485: out <= 16'h054C;    16'd47486: out <= 16'hF9FC;    16'd47487: out <= 16'h0518;
    16'd47488: out <= 16'hFF20;    16'd47489: out <= 16'hF9BA;    16'd47490: out <= 16'hFF54;    16'd47491: out <= 16'hFBC3;
    16'd47492: out <= 16'h00DD;    16'd47493: out <= 16'hFEB1;    16'd47494: out <= 16'hFE48;    16'd47495: out <= 16'h0448;
    16'd47496: out <= 16'h0502;    16'd47497: out <= 16'hFC51;    16'd47498: out <= 16'h00B6;    16'd47499: out <= 16'hFF0C;
    16'd47500: out <= 16'h0187;    16'd47501: out <= 16'h01B1;    16'd47502: out <= 16'hFE43;    16'd47503: out <= 16'hFE72;
    16'd47504: out <= 16'h00A2;    16'd47505: out <= 16'h0068;    16'd47506: out <= 16'hFCE2;    16'd47507: out <= 16'hFFFA;
    16'd47508: out <= 16'hFFC6;    16'd47509: out <= 16'hFDE4;    16'd47510: out <= 16'h000E;    16'd47511: out <= 16'hFF1C;
    16'd47512: out <= 16'hFC06;    16'd47513: out <= 16'hFB1D;    16'd47514: out <= 16'h014D;    16'd47515: out <= 16'hFE66;
    16'd47516: out <= 16'h0032;    16'd47517: out <= 16'h0321;    16'd47518: out <= 16'h005E;    16'd47519: out <= 16'h03AA;
    16'd47520: out <= 16'h03A3;    16'd47521: out <= 16'h0188;    16'd47522: out <= 16'h0AF4;    16'd47523: out <= 16'h0D32;
    16'd47524: out <= 16'h04F9;    16'd47525: out <= 16'h01D4;    16'd47526: out <= 16'h0636;    16'd47527: out <= 16'h00B3;
    16'd47528: out <= 16'h0A39;    16'd47529: out <= 16'h04F2;    16'd47530: out <= 16'hFCEE;    16'd47531: out <= 16'h0746;
    16'd47532: out <= 16'h039A;    16'd47533: out <= 16'h0535;    16'd47534: out <= 16'hFF27;    16'd47535: out <= 16'h046E;
    16'd47536: out <= 16'h00E0;    16'd47537: out <= 16'h01D6;    16'd47538: out <= 16'h0774;    16'd47539: out <= 16'h0BF6;
    16'd47540: out <= 16'h052F;    16'd47541: out <= 16'h0677;    16'd47542: out <= 16'h0581;    16'd47543: out <= 16'h0447;
    16'd47544: out <= 16'hFB03;    16'd47545: out <= 16'hFF23;    16'd47546: out <= 16'h0892;    16'd47547: out <= 16'h0264;
    16'd47548: out <= 16'h0134;    16'd47549: out <= 16'h05C9;    16'd47550: out <= 16'h0107;    16'd47551: out <= 16'h0BB0;
    16'd47552: out <= 16'h02F4;    16'd47553: out <= 16'h08DC;    16'd47554: out <= 16'h06C5;    16'd47555: out <= 16'hFC70;
    16'd47556: out <= 16'h04B6;    16'd47557: out <= 16'h0AFA;    16'd47558: out <= 16'h0564;    16'd47559: out <= 16'h03B1;
    16'd47560: out <= 16'h005C;    16'd47561: out <= 16'hF686;    16'd47562: out <= 16'hFB09;    16'd47563: out <= 16'h021A;
    16'd47564: out <= 16'h064A;    16'd47565: out <= 16'h009E;    16'd47566: out <= 16'hFD13;    16'd47567: out <= 16'hF7EB;
    16'd47568: out <= 16'hFECB;    16'd47569: out <= 16'hFC88;    16'd47570: out <= 16'h012F;    16'd47571: out <= 16'h0390;
    16'd47572: out <= 16'hFE91;    16'd47573: out <= 16'hF87B;    16'd47574: out <= 16'h050E;    16'd47575: out <= 16'h0100;
    16'd47576: out <= 16'h002F;    16'd47577: out <= 16'hF8F8;    16'd47578: out <= 16'h080E;    16'd47579: out <= 16'hFD3D;
    16'd47580: out <= 16'h0A9F;    16'd47581: out <= 16'hFFBE;    16'd47582: out <= 16'h0063;    16'd47583: out <= 16'h0068;
    16'd47584: out <= 16'hF787;    16'd47585: out <= 16'h0384;    16'd47586: out <= 16'hFE3A;    16'd47587: out <= 16'h0061;
    16'd47588: out <= 16'hF8AA;    16'd47589: out <= 16'h0245;    16'd47590: out <= 16'h0165;    16'd47591: out <= 16'h02CE;
    16'd47592: out <= 16'h0663;    16'd47593: out <= 16'hFFFA;    16'd47594: out <= 16'h0561;    16'd47595: out <= 16'h017B;
    16'd47596: out <= 16'h043E;    16'd47597: out <= 16'h02E2;    16'd47598: out <= 16'h0359;    16'd47599: out <= 16'hFF2B;
    16'd47600: out <= 16'hFD7E;    16'd47601: out <= 16'hFE9E;    16'd47602: out <= 16'h0398;    16'd47603: out <= 16'hFE9D;
    16'd47604: out <= 16'h0303;    16'd47605: out <= 16'h040B;    16'd47606: out <= 16'hFD87;    16'd47607: out <= 16'hFDE5;
    16'd47608: out <= 16'hFD54;    16'd47609: out <= 16'hFE20;    16'd47610: out <= 16'hF9D7;    16'd47611: out <= 16'hFE45;
    16'd47612: out <= 16'h01BE;    16'd47613: out <= 16'h00BF;    16'd47614: out <= 16'hFBC9;    16'd47615: out <= 16'h002B;
    16'd47616: out <= 16'h0128;    16'd47617: out <= 16'hFBCA;    16'd47618: out <= 16'hF9EF;    16'd47619: out <= 16'h04E5;
    16'd47620: out <= 16'h0045;    16'd47621: out <= 16'hFFF3;    16'd47622: out <= 16'hF9B2;    16'd47623: out <= 16'h017D;
    16'd47624: out <= 16'hFF75;    16'd47625: out <= 16'hFC1E;    16'd47626: out <= 16'hFED1;    16'd47627: out <= 16'h08D7;
    16'd47628: out <= 16'hFFD5;    16'd47629: out <= 16'hFB19;    16'd47630: out <= 16'hFCDF;    16'd47631: out <= 16'hFF18;
    16'd47632: out <= 16'h0276;    16'd47633: out <= 16'hF965;    16'd47634: out <= 16'h0051;    16'd47635: out <= 16'h02A4;
    16'd47636: out <= 16'hFF8A;    16'd47637: out <= 16'h05B9;    16'd47638: out <= 16'hFEA9;    16'd47639: out <= 16'h02CC;
    16'd47640: out <= 16'hFF9E;    16'd47641: out <= 16'hF867;    16'd47642: out <= 16'hF7BF;    16'd47643: out <= 16'hFBD0;
    16'd47644: out <= 16'hFD14;    16'd47645: out <= 16'hFAC2;    16'd47646: out <= 16'h0338;    16'd47647: out <= 16'h0030;
    16'd47648: out <= 16'hFF1D;    16'd47649: out <= 16'hFD51;    16'd47650: out <= 16'h01D8;    16'd47651: out <= 16'h0250;
    16'd47652: out <= 16'h0127;    16'd47653: out <= 16'hFE28;    16'd47654: out <= 16'h02F9;    16'd47655: out <= 16'h05CB;
    16'd47656: out <= 16'h018C;    16'd47657: out <= 16'h09B3;    16'd47658: out <= 16'h04DD;    16'd47659: out <= 16'h1022;
    16'd47660: out <= 16'h044B;    16'd47661: out <= 16'hFD68;    16'd47662: out <= 16'hF766;    16'd47663: out <= 16'h06A1;
    16'd47664: out <= 16'h0178;    16'd47665: out <= 16'h0691;    16'd47666: out <= 16'h0A5A;    16'd47667: out <= 16'h0548;
    16'd47668: out <= 16'h0215;    16'd47669: out <= 16'h0329;    16'd47670: out <= 16'h00CB;    16'd47671: out <= 16'h02D1;
    16'd47672: out <= 16'h09CB;    16'd47673: out <= 16'h0227;    16'd47674: out <= 16'h05F7;    16'd47675: out <= 16'h00F4;
    16'd47676: out <= 16'hFED9;    16'd47677: out <= 16'h0C00;    16'd47678: out <= 16'h075F;    16'd47679: out <= 16'h03C0;
    16'd47680: out <= 16'h0223;    16'd47681: out <= 16'h03EC;    16'd47682: out <= 16'h0A35;    16'd47683: out <= 16'h07DB;
    16'd47684: out <= 16'h04C5;    16'd47685: out <= 16'h04AE;    16'd47686: out <= 16'h0404;    16'd47687: out <= 16'h028E;
    16'd47688: out <= 16'hFE85;    16'd47689: out <= 16'h0579;    16'd47690: out <= 16'h0B27;    16'd47691: out <= 16'hF9DB;
    16'd47692: out <= 16'hFDA4;    16'd47693: out <= 16'h0614;    16'd47694: out <= 16'h0422;    16'd47695: out <= 16'h07D4;
    16'd47696: out <= 16'h0026;    16'd47697: out <= 16'h048C;    16'd47698: out <= 16'h02AE;    16'd47699: out <= 16'h0126;
    16'd47700: out <= 16'h0142;    16'd47701: out <= 16'h0262;    16'd47702: out <= 16'hFE3F;    16'd47703: out <= 16'h055C;
    16'd47704: out <= 16'hFD4C;    16'd47705: out <= 16'h01A8;    16'd47706: out <= 16'h03CE;    16'd47707: out <= 16'h01CA;
    16'd47708: out <= 16'h0159;    16'd47709: out <= 16'h03B0;    16'd47710: out <= 16'hF7A6;    16'd47711: out <= 16'h032E;
    16'd47712: out <= 16'h062F;    16'd47713: out <= 16'h0434;    16'd47714: out <= 16'h0458;    16'd47715: out <= 16'hFD95;
    16'd47716: out <= 16'h0237;    16'd47717: out <= 16'h0C8C;    16'd47718: out <= 16'h0114;    16'd47719: out <= 16'h03E9;
    16'd47720: out <= 16'hFC0A;    16'd47721: out <= 16'h049F;    16'd47722: out <= 16'hF7D0;    16'd47723: out <= 16'h00CE;
    16'd47724: out <= 16'hFD83;    16'd47725: out <= 16'hFD8F;    16'd47726: out <= 16'hF95A;    16'd47727: out <= 16'hFFF5;
    16'd47728: out <= 16'h089A;    16'd47729: out <= 16'hFDF0;    16'd47730: out <= 16'hFD21;    16'd47731: out <= 16'hFF40;
    16'd47732: out <= 16'hFC6E;    16'd47733: out <= 16'h0027;    16'd47734: out <= 16'hFCB9;    16'd47735: out <= 16'hFC46;
    16'd47736: out <= 16'h0522;    16'd47737: out <= 16'hFFFE;    16'd47738: out <= 16'h017A;    16'd47739: out <= 16'h010B;
    16'd47740: out <= 16'h04BD;    16'd47741: out <= 16'hFC5B;    16'd47742: out <= 16'h048D;    16'd47743: out <= 16'hFE7F;
    16'd47744: out <= 16'hFAD1;    16'd47745: out <= 16'h00A3;    16'd47746: out <= 16'hFD2B;    16'd47747: out <= 16'h00E4;
    16'd47748: out <= 16'hFC80;    16'd47749: out <= 16'hFE00;    16'd47750: out <= 16'hFAB6;    16'd47751: out <= 16'hFB25;
    16'd47752: out <= 16'h090C;    16'd47753: out <= 16'h04DF;    16'd47754: out <= 16'h0225;    16'd47755: out <= 16'h0475;
    16'd47756: out <= 16'h00C1;    16'd47757: out <= 16'h0420;    16'd47758: out <= 16'hF813;    16'd47759: out <= 16'hFCDD;
    16'd47760: out <= 16'hFF06;    16'd47761: out <= 16'h0499;    16'd47762: out <= 16'hFB6A;    16'd47763: out <= 16'h0A7C;
    16'd47764: out <= 16'h039B;    16'd47765: out <= 16'h01E8;    16'd47766: out <= 16'hFBD5;    16'd47767: out <= 16'hF783;
    16'd47768: out <= 16'h017D;    16'd47769: out <= 16'h04DD;    16'd47770: out <= 16'hFBD4;    16'd47771: out <= 16'hFC11;
    16'd47772: out <= 16'h04DA;    16'd47773: out <= 16'h0015;    16'd47774: out <= 16'h0038;    16'd47775: out <= 16'h0018;
    16'd47776: out <= 16'h04E1;    16'd47777: out <= 16'h073D;    16'd47778: out <= 16'h050E;    16'd47779: out <= 16'h0752;
    16'd47780: out <= 16'h091A;    16'd47781: out <= 16'h0199;    16'd47782: out <= 16'h0416;    16'd47783: out <= 16'h0038;
    16'd47784: out <= 16'hFF82;    16'd47785: out <= 16'h0266;    16'd47786: out <= 16'hFFEC;    16'd47787: out <= 16'h019C;
    16'd47788: out <= 16'h04F1;    16'd47789: out <= 16'h01BE;    16'd47790: out <= 16'h0023;    16'd47791: out <= 16'h031B;
    16'd47792: out <= 16'h06BF;    16'd47793: out <= 16'hFEA2;    16'd47794: out <= 16'h06BC;    16'd47795: out <= 16'h092C;
    16'd47796: out <= 16'h081F;    16'd47797: out <= 16'h0249;    16'd47798: out <= 16'hFC27;    16'd47799: out <= 16'h03EA;
    16'd47800: out <= 16'h0547;    16'd47801: out <= 16'h0073;    16'd47802: out <= 16'h010D;    16'd47803: out <= 16'hFFEF;
    16'd47804: out <= 16'h0547;    16'd47805: out <= 16'hFBD7;    16'd47806: out <= 16'h04C0;    16'd47807: out <= 16'h09C0;
    16'd47808: out <= 16'h04E6;    16'd47809: out <= 16'h0494;    16'd47810: out <= 16'h0959;    16'd47811: out <= 16'hFE9A;
    16'd47812: out <= 16'hFE73;    16'd47813: out <= 16'h02EB;    16'd47814: out <= 16'h09B4;    16'd47815: out <= 16'h0535;
    16'd47816: out <= 16'hFDCC;    16'd47817: out <= 16'hF8E5;    16'd47818: out <= 16'hFD41;    16'd47819: out <= 16'h0515;
    16'd47820: out <= 16'h0707;    16'd47821: out <= 16'h03E1;    16'd47822: out <= 16'hFB4B;    16'd47823: out <= 16'h0863;
    16'd47824: out <= 16'h009C;    16'd47825: out <= 16'h0590;    16'd47826: out <= 16'h04F6;    16'd47827: out <= 16'hFD21;
    16'd47828: out <= 16'hFC22;    16'd47829: out <= 16'h06F6;    16'd47830: out <= 16'hFEE9;    16'd47831: out <= 16'h015B;
    16'd47832: out <= 16'hF975;    16'd47833: out <= 16'h02A1;    16'd47834: out <= 16'hFFDC;    16'd47835: out <= 16'hFD2A;
    16'd47836: out <= 16'hFDE4;    16'd47837: out <= 16'h01B8;    16'd47838: out <= 16'h01CE;    16'd47839: out <= 16'hFDA3;
    16'd47840: out <= 16'hFEA8;    16'd47841: out <= 16'hFBD5;    16'd47842: out <= 16'hF936;    16'd47843: out <= 16'hFD5E;
    16'd47844: out <= 16'hFF08;    16'd47845: out <= 16'h0166;    16'd47846: out <= 16'hFD19;    16'd47847: out <= 16'hFFA9;
    16'd47848: out <= 16'h025D;    16'd47849: out <= 16'hFB94;    16'd47850: out <= 16'h02C8;    16'd47851: out <= 16'h0125;
    16'd47852: out <= 16'h057C;    16'd47853: out <= 16'h04BD;    16'd47854: out <= 16'h0021;    16'd47855: out <= 16'h04E8;
    16'd47856: out <= 16'hFE67;    16'd47857: out <= 16'hF9FD;    16'd47858: out <= 16'hFB39;    16'd47859: out <= 16'h0322;
    16'd47860: out <= 16'hFF69;    16'd47861: out <= 16'h068C;    16'd47862: out <= 16'h053A;    16'd47863: out <= 16'h0893;
    16'd47864: out <= 16'h026B;    16'd47865: out <= 16'hF7AE;    16'd47866: out <= 16'hFC31;    16'd47867: out <= 16'hFEC8;
    16'd47868: out <= 16'h071E;    16'd47869: out <= 16'h0137;    16'd47870: out <= 16'hFE99;    16'd47871: out <= 16'h0202;
    16'd47872: out <= 16'h0006;    16'd47873: out <= 16'h02D7;    16'd47874: out <= 16'hFE5C;    16'd47875: out <= 16'h020A;
    16'd47876: out <= 16'hFCFE;    16'd47877: out <= 16'hFE35;    16'd47878: out <= 16'hFDAD;    16'd47879: out <= 16'h074A;
    16'd47880: out <= 16'hFE8E;    16'd47881: out <= 16'h020F;    16'd47882: out <= 16'h0456;    16'd47883: out <= 16'h015D;
    16'd47884: out <= 16'h049A;    16'd47885: out <= 16'h01FB;    16'd47886: out <= 16'hFA9D;    16'd47887: out <= 16'h0412;
    16'd47888: out <= 16'hFCAF;    16'd47889: out <= 16'hFBDA;    16'd47890: out <= 16'hFEB8;    16'd47891: out <= 16'hF967;
    16'd47892: out <= 16'h0075;    16'd47893: out <= 16'hFBE7;    16'd47894: out <= 16'hF905;    16'd47895: out <= 16'hFF8F;
    16'd47896: out <= 16'h0310;    16'd47897: out <= 16'h06DC;    16'd47898: out <= 16'hF9B1;    16'd47899: out <= 16'hFDE9;
    16'd47900: out <= 16'hFB8E;    16'd47901: out <= 16'h00E2;    16'd47902: out <= 16'h0513;    16'd47903: out <= 16'hFAA5;
    16'd47904: out <= 16'hFBE7;    16'd47905: out <= 16'h0111;    16'd47906: out <= 16'hFF5D;    16'd47907: out <= 16'h05BC;
    16'd47908: out <= 16'h06AA;    16'd47909: out <= 16'h0370;    16'd47910: out <= 16'h0451;    16'd47911: out <= 16'hFFBD;
    16'd47912: out <= 16'h0D33;    16'd47913: out <= 16'h0879;    16'd47914: out <= 16'hFEB4;    16'd47915: out <= 16'h03FE;
    16'd47916: out <= 16'h0475;    16'd47917: out <= 16'h04A0;    16'd47918: out <= 16'h0400;    16'd47919: out <= 16'h0021;
    16'd47920: out <= 16'h025C;    16'd47921: out <= 16'h05AC;    16'd47922: out <= 16'h08FA;    16'd47923: out <= 16'h0620;
    16'd47924: out <= 16'h0508;    16'd47925: out <= 16'h0645;    16'd47926: out <= 16'h05CB;    16'd47927: out <= 16'h061A;
    16'd47928: out <= 16'h03A2;    16'd47929: out <= 16'h0893;    16'd47930: out <= 16'hFD86;    16'd47931: out <= 16'h07D8;
    16'd47932: out <= 16'hFEC2;    16'd47933: out <= 16'h0460;    16'd47934: out <= 16'h0470;    16'd47935: out <= 16'hFE48;
    16'd47936: out <= 16'h078C;    16'd47937: out <= 16'h0681;    16'd47938: out <= 16'h05B2;    16'd47939: out <= 16'h047D;
    16'd47940: out <= 16'h0164;    16'd47941: out <= 16'hFEDF;    16'd47942: out <= 16'hFEF6;    16'd47943: out <= 16'h041A;
    16'd47944: out <= 16'h08F5;    16'd47945: out <= 16'h06BC;    16'd47946: out <= 16'h0B2F;    16'd47947: out <= 16'h031F;
    16'd47948: out <= 16'h064C;    16'd47949: out <= 16'h0B0C;    16'd47950: out <= 16'h068F;    16'd47951: out <= 16'h05C2;
    16'd47952: out <= 16'h0387;    16'd47953: out <= 16'h0175;    16'd47954: out <= 16'h0682;    16'd47955: out <= 16'h0047;
    16'd47956: out <= 16'h0820;    16'd47957: out <= 16'h0427;    16'd47958: out <= 16'h0750;    16'd47959: out <= 16'h01BD;
    16'd47960: out <= 16'h02D7;    16'd47961: out <= 16'h005E;    16'd47962: out <= 16'h0686;    16'd47963: out <= 16'h016F;
    16'd47964: out <= 16'h026B;    16'd47965: out <= 16'h02CB;    16'd47966: out <= 16'h02D0;    16'd47967: out <= 16'h0337;
    16'd47968: out <= 16'h0198;    16'd47969: out <= 16'h010B;    16'd47970: out <= 16'h070F;    16'd47971: out <= 16'h05A7;
    16'd47972: out <= 16'h0219;    16'd47973: out <= 16'h057A;    16'd47974: out <= 16'h0664;    16'd47975: out <= 16'h05F7;
    16'd47976: out <= 16'h060F;    16'd47977: out <= 16'h06BA;    16'd47978: out <= 16'hFF67;    16'd47979: out <= 16'h0920;
    16'd47980: out <= 16'h01FF;    16'd47981: out <= 16'hFE5B;    16'd47982: out <= 16'h0265;    16'd47983: out <= 16'h075D;
    16'd47984: out <= 16'hFF7F;    16'd47985: out <= 16'hFB3A;    16'd47986: out <= 16'hF57D;    16'd47987: out <= 16'h0015;
    16'd47988: out <= 16'h0370;    16'd47989: out <= 16'hFA39;    16'd47990: out <= 16'hF99D;    16'd47991: out <= 16'hFF0A;
    16'd47992: out <= 16'h072D;    16'd47993: out <= 16'hFFF1;    16'd47994: out <= 16'hFC7E;    16'd47995: out <= 16'h009F;
    16'd47996: out <= 16'h00D4;    16'd47997: out <= 16'h0215;    16'd47998: out <= 16'h04F3;    16'd47999: out <= 16'hFCFA;
    16'd48000: out <= 16'h0079;    16'd48001: out <= 16'h0371;    16'd48002: out <= 16'h0433;    16'd48003: out <= 16'hFE7C;
    16'd48004: out <= 16'h0191;    16'd48005: out <= 16'h0008;    16'd48006: out <= 16'h04C3;    16'd48007: out <= 16'hFF0F;
    16'd48008: out <= 16'h01DD;    16'd48009: out <= 16'hFD37;    16'd48010: out <= 16'h0333;    16'd48011: out <= 16'h0310;
    16'd48012: out <= 16'h0213;    16'd48013: out <= 16'h0151;    16'd48014: out <= 16'hFA1B;    16'd48015: out <= 16'hFD6D;
    16'd48016: out <= 16'hFDA2;    16'd48017: out <= 16'h083C;    16'd48018: out <= 16'h03E7;    16'd48019: out <= 16'hFC57;
    16'd48020: out <= 16'h0390;    16'd48021: out <= 16'h01D7;    16'd48022: out <= 16'h026F;    16'd48023: out <= 16'h0397;
    16'd48024: out <= 16'h016B;    16'd48025: out <= 16'h0A1C;    16'd48026: out <= 16'h0360;    16'd48027: out <= 16'h0079;
    16'd48028: out <= 16'h039C;    16'd48029: out <= 16'h0213;    16'd48030: out <= 16'h093E;    16'd48031: out <= 16'h0735;
    16'd48032: out <= 16'h0670;    16'd48033: out <= 16'h073A;    16'd48034: out <= 16'h031A;    16'd48035: out <= 16'h04E0;
    16'd48036: out <= 16'hFE62;    16'd48037: out <= 16'h019B;    16'd48038: out <= 16'h02EE;    16'd48039: out <= 16'h0787;
    16'd48040: out <= 16'h01C9;    16'd48041: out <= 16'h091F;    16'd48042: out <= 16'h01F5;    16'd48043: out <= 16'h04A2;
    16'd48044: out <= 16'h0632;    16'd48045: out <= 16'h03CA;    16'd48046: out <= 16'hFE7C;    16'd48047: out <= 16'h077F;
    16'd48048: out <= 16'h0579;    16'd48049: out <= 16'h0318;    16'd48050: out <= 16'h04A3;    16'd48051: out <= 16'h0448;
    16'd48052: out <= 16'h016A;    16'd48053: out <= 16'h0689;    16'd48054: out <= 16'h0499;    16'd48055: out <= 16'h0357;
    16'd48056: out <= 16'h0451;    16'd48057: out <= 16'h0011;    16'd48058: out <= 16'h0754;    16'd48059: out <= 16'hFCCA;
    16'd48060: out <= 16'hFEE8;    16'd48061: out <= 16'h02A3;    16'd48062: out <= 16'h0316;    16'd48063: out <= 16'h057C;
    16'd48064: out <= 16'h049A;    16'd48065: out <= 16'h01EC;    16'd48066: out <= 16'h059E;    16'd48067: out <= 16'h001A;
    16'd48068: out <= 16'hFFC4;    16'd48069: out <= 16'hF6C6;    16'd48070: out <= 16'h012E;    16'd48071: out <= 16'h0263;
    16'd48072: out <= 16'hFB7A;    16'd48073: out <= 16'h0269;    16'd48074: out <= 16'h00A8;    16'd48075: out <= 16'hFDCF;
    16'd48076: out <= 16'h05DF;    16'd48077: out <= 16'hFAE0;    16'd48078: out <= 16'h070A;    16'd48079: out <= 16'hFC22;
    16'd48080: out <= 16'h0484;    16'd48081: out <= 16'h0424;    16'd48082: out <= 16'h030E;    16'd48083: out <= 16'h0288;
    16'd48084: out <= 16'hFF72;    16'd48085: out <= 16'hFCBA;    16'd48086: out <= 16'hFFAD;    16'd48087: out <= 16'h019E;
    16'd48088: out <= 16'hF911;    16'd48089: out <= 16'hFBC9;    16'd48090: out <= 16'hFF38;    16'd48091: out <= 16'h0394;
    16'd48092: out <= 16'h0264;    16'd48093: out <= 16'hFBFC;    16'd48094: out <= 16'h00E0;    16'd48095: out <= 16'hFED8;
    16'd48096: out <= 16'hFA11;    16'd48097: out <= 16'hFAF8;    16'd48098: out <= 16'hFC7F;    16'd48099: out <= 16'hFB62;
    16'd48100: out <= 16'h018D;    16'd48101: out <= 16'h027D;    16'd48102: out <= 16'h0491;    16'd48103: out <= 16'hFF20;
    16'd48104: out <= 16'hFD58;    16'd48105: out <= 16'h00EA;    16'd48106: out <= 16'h0484;    16'd48107: out <= 16'hFE03;
    16'd48108: out <= 16'hFD1A;    16'd48109: out <= 16'h0002;    16'd48110: out <= 16'hF981;    16'd48111: out <= 16'h0471;
    16'd48112: out <= 16'h0217;    16'd48113: out <= 16'h0250;    16'd48114: out <= 16'hF940;    16'd48115: out <= 16'hF9D9;
    16'd48116: out <= 16'hFBCC;    16'd48117: out <= 16'h03DC;    16'd48118: out <= 16'h03FD;    16'd48119: out <= 16'h00C7;
    16'd48120: out <= 16'hFAD4;    16'd48121: out <= 16'hFB46;    16'd48122: out <= 16'hFF47;    16'd48123: out <= 16'hFFA6;
    16'd48124: out <= 16'hFA1B;    16'd48125: out <= 16'h026C;    16'd48126: out <= 16'hFF2F;    16'd48127: out <= 16'hFF9C;
    16'd48128: out <= 16'h06CF;    16'd48129: out <= 16'hFEB4;    16'd48130: out <= 16'h02C0;    16'd48131: out <= 16'hF9C4;
    16'd48132: out <= 16'h0069;    16'd48133: out <= 16'hFF6F;    16'd48134: out <= 16'h01F9;    16'd48135: out <= 16'hFCDB;
    16'd48136: out <= 16'hFCB5;    16'd48137: out <= 16'hFEAA;    16'd48138: out <= 16'h04C9;    16'd48139: out <= 16'h0221;
    16'd48140: out <= 16'hFF83;    16'd48141: out <= 16'h01F7;    16'd48142: out <= 16'h06EA;    16'd48143: out <= 16'hFD80;
    16'd48144: out <= 16'h029D;    16'd48145: out <= 16'h03E8;    16'd48146: out <= 16'h051B;    16'd48147: out <= 16'h01EF;
    16'd48148: out <= 16'h0264;    16'd48149: out <= 16'hFA13;    16'd48150: out <= 16'h00DC;    16'd48151: out <= 16'h0286;
    16'd48152: out <= 16'hF6A3;    16'd48153: out <= 16'h0429;    16'd48154: out <= 16'hFFF6;    16'd48155: out <= 16'hFE3C;
    16'd48156: out <= 16'h01C2;    16'd48157: out <= 16'h03CB;    16'd48158: out <= 16'hFE92;    16'd48159: out <= 16'h0381;
    16'd48160: out <= 16'h01C7;    16'd48161: out <= 16'hFA46;    16'd48162: out <= 16'h01A4;    16'd48163: out <= 16'h0111;
    16'd48164: out <= 16'hFF1A;    16'd48165: out <= 16'hFB86;    16'd48166: out <= 16'hFBDE;    16'd48167: out <= 16'h018C;
    16'd48168: out <= 16'h01BB;    16'd48169: out <= 16'h04D5;    16'd48170: out <= 16'h03A6;    16'd48171: out <= 16'h0332;
    16'd48172: out <= 16'h031A;    16'd48173: out <= 16'h0279;    16'd48174: out <= 16'h01FA;    16'd48175: out <= 16'h0293;
    16'd48176: out <= 16'h00A5;    16'd48177: out <= 16'h03D4;    16'd48178: out <= 16'h074B;    16'd48179: out <= 16'h0415;
    16'd48180: out <= 16'h04EB;    16'd48181: out <= 16'hFD87;    16'd48182: out <= 16'h0AA5;    16'd48183: out <= 16'h0238;
    16'd48184: out <= 16'h0475;    16'd48185: out <= 16'h0021;    16'd48186: out <= 16'h0768;    16'd48187: out <= 16'h0619;
    16'd48188: out <= 16'h0107;    16'd48189: out <= 16'hFBF9;    16'd48190: out <= 16'hFF61;    16'd48191: out <= 16'hFC4D;
    16'd48192: out <= 16'hFBFE;    16'd48193: out <= 16'h07CF;    16'd48194: out <= 16'h0308;    16'd48195: out <= 16'h03EC;
    16'd48196: out <= 16'h0478;    16'd48197: out <= 16'h0118;    16'd48198: out <= 16'h05C5;    16'd48199: out <= 16'h0871;
    16'd48200: out <= 16'h03D5;    16'd48201: out <= 16'hFDE6;    16'd48202: out <= 16'h044A;    16'd48203: out <= 16'hFFF9;
    16'd48204: out <= 16'h0775;    16'd48205: out <= 16'h0037;    16'd48206: out <= 16'h0551;    16'd48207: out <= 16'h0A96;
    16'd48208: out <= 16'h07D7;    16'd48209: out <= 16'h0377;    16'd48210: out <= 16'h0196;    16'd48211: out <= 16'hFF4C;
    16'd48212: out <= 16'h0241;    16'd48213: out <= 16'h06D1;    16'd48214: out <= 16'h0237;    16'd48215: out <= 16'h0082;
    16'd48216: out <= 16'h02A7;    16'd48217: out <= 16'h04F7;    16'd48218: out <= 16'h09AE;    16'd48219: out <= 16'hFF53;
    16'd48220: out <= 16'h0089;    16'd48221: out <= 16'h04EB;    16'd48222: out <= 16'hFF52;    16'd48223: out <= 16'h0078;
    16'd48224: out <= 16'hFC60;    16'd48225: out <= 16'h02CD;    16'd48226: out <= 16'h01BA;    16'd48227: out <= 16'h05CE;
    16'd48228: out <= 16'h0AAE;    16'd48229: out <= 16'h0213;    16'd48230: out <= 16'h0237;    16'd48231: out <= 16'hFD52;
    16'd48232: out <= 16'h0105;    16'd48233: out <= 16'h03FE;    16'd48234: out <= 16'h009B;    16'd48235: out <= 16'h021B;
    16'd48236: out <= 16'h0097;    16'd48237: out <= 16'h03F1;    16'd48238: out <= 16'hFDCD;    16'd48239: out <= 16'h010D;
    16'd48240: out <= 16'hFDEB;    16'd48241: out <= 16'h0A8F;    16'd48242: out <= 16'h013D;    16'd48243: out <= 16'h094D;
    16'd48244: out <= 16'h00E2;    16'd48245: out <= 16'h00C3;    16'd48246: out <= 16'h03D6;    16'd48247: out <= 16'hFFCF;
    16'd48248: out <= 16'h0A74;    16'd48249: out <= 16'hFD72;    16'd48250: out <= 16'h02FB;    16'd48251: out <= 16'h0186;
    16'd48252: out <= 16'h00CF;    16'd48253: out <= 16'h015E;    16'd48254: out <= 16'h04DC;    16'd48255: out <= 16'h05C1;
    16'd48256: out <= 16'h0301;    16'd48257: out <= 16'h057A;    16'd48258: out <= 16'h02D3;    16'd48259: out <= 16'h074A;
    16'd48260: out <= 16'hFD82;    16'd48261: out <= 16'hFF9F;    16'd48262: out <= 16'hFFC2;    16'd48263: out <= 16'h050F;
    16'd48264: out <= 16'h0382;    16'd48265: out <= 16'h020C;    16'd48266: out <= 16'h00B8;    16'd48267: out <= 16'h032D;
    16'd48268: out <= 16'h0097;    16'd48269: out <= 16'hFF2E;    16'd48270: out <= 16'hFE7D;    16'd48271: out <= 16'h0889;
    16'd48272: out <= 16'h07A9;    16'd48273: out <= 16'h06A0;    16'd48274: out <= 16'hFAA5;    16'd48275: out <= 16'h06F7;
    16'd48276: out <= 16'h0011;    16'd48277: out <= 16'hFC36;    16'd48278: out <= 16'h01DD;    16'd48279: out <= 16'hFF8B;
    16'd48280: out <= 16'hFDD6;    16'd48281: out <= 16'h03AF;    16'd48282: out <= 16'hF92E;    16'd48283: out <= 16'hFC02;
    16'd48284: out <= 16'h0A4D;    16'd48285: out <= 16'h01C2;    16'd48286: out <= 16'h0737;    16'd48287: out <= 16'hFF90;
    16'd48288: out <= 16'h07FE;    16'd48289: out <= 16'hFF39;    16'd48290: out <= 16'h02DD;    16'd48291: out <= 16'h07CF;
    16'd48292: out <= 16'h028D;    16'd48293: out <= 16'h0512;    16'd48294: out <= 16'h0413;    16'd48295: out <= 16'h0166;
    16'd48296: out <= 16'h03F3;    16'd48297: out <= 16'h0538;    16'd48298: out <= 16'h04AC;    16'd48299: out <= 16'h075B;
    16'd48300: out <= 16'h006D;    16'd48301: out <= 16'h065D;    16'd48302: out <= 16'h040E;    16'd48303: out <= 16'h03FC;
    16'd48304: out <= 16'hFC34;    16'd48305: out <= 16'h0319;    16'd48306: out <= 16'h06F2;    16'd48307: out <= 16'h0890;
    16'd48308: out <= 16'h0393;    16'd48309: out <= 16'hFD4A;    16'd48310: out <= 16'hFEBC;    16'd48311: out <= 16'h0884;
    16'd48312: out <= 16'h058D;    16'd48313: out <= 16'h08D9;    16'd48314: out <= 16'h05A6;    16'd48315: out <= 16'hF8D0;
    16'd48316: out <= 16'h028C;    16'd48317: out <= 16'h0073;    16'd48318: out <= 16'h040C;    16'd48319: out <= 16'h014A;
    16'd48320: out <= 16'h052D;    16'd48321: out <= 16'h00C2;    16'd48322: out <= 16'h0710;    16'd48323: out <= 16'h0006;
    16'd48324: out <= 16'h0536;    16'd48325: out <= 16'h02D2;    16'd48326: out <= 16'h0384;    16'd48327: out <= 16'h02D4;
    16'd48328: out <= 16'h0421;    16'd48329: out <= 16'hF9FE;    16'd48330: out <= 16'h00BC;    16'd48331: out <= 16'h04A6;
    16'd48332: out <= 16'hFEFF;    16'd48333: out <= 16'h004B;    16'd48334: out <= 16'hFB69;    16'd48335: out <= 16'h020E;
    16'd48336: out <= 16'h0C1C;    16'd48337: out <= 16'h0523;    16'd48338: out <= 16'hFF27;    16'd48339: out <= 16'hFD11;
    16'd48340: out <= 16'h03FC;    16'd48341: out <= 16'h0436;    16'd48342: out <= 16'h0176;    16'd48343: out <= 16'h05A3;
    16'd48344: out <= 16'h021F;    16'd48345: out <= 16'hFCD0;    16'd48346: out <= 16'hFE8D;    16'd48347: out <= 16'h0305;
    16'd48348: out <= 16'hFFBC;    16'd48349: out <= 16'hFD2C;    16'd48350: out <= 16'h0040;    16'd48351: out <= 16'hFC3A;
    16'd48352: out <= 16'hFFAB;    16'd48353: out <= 16'hFB2D;    16'd48354: out <= 16'hFF3A;    16'd48355: out <= 16'h0133;
    16'd48356: out <= 16'hFC63;    16'd48357: out <= 16'hF83D;    16'd48358: out <= 16'h02A4;    16'd48359: out <= 16'hF833;
    16'd48360: out <= 16'h0161;    16'd48361: out <= 16'hF54E;    16'd48362: out <= 16'h0695;    16'd48363: out <= 16'hFDE6;
    16'd48364: out <= 16'h07A6;    16'd48365: out <= 16'h0124;    16'd48366: out <= 16'h011A;    16'd48367: out <= 16'hFD52;
    16'd48368: out <= 16'hFCBD;    16'd48369: out <= 16'hFF4A;    16'd48370: out <= 16'h00B7;    16'd48371: out <= 16'hF89D;
    16'd48372: out <= 16'hF9DA;    16'd48373: out <= 16'hFF7A;    16'd48374: out <= 16'hFDAE;    16'd48375: out <= 16'h0005;
    16'd48376: out <= 16'hF87B;    16'd48377: out <= 16'h01CB;    16'd48378: out <= 16'h05DE;    16'd48379: out <= 16'h0068;
    16'd48380: out <= 16'h036E;    16'd48381: out <= 16'hFEFF;    16'd48382: out <= 16'hFFCA;    16'd48383: out <= 16'h0351;
    16'd48384: out <= 16'hFCF7;    16'd48385: out <= 16'h01B8;    16'd48386: out <= 16'h0042;    16'd48387: out <= 16'h023D;
    16'd48388: out <= 16'h001E;    16'd48389: out <= 16'hF88D;    16'd48390: out <= 16'h0634;    16'd48391: out <= 16'h03E3;
    16'd48392: out <= 16'h0305;    16'd48393: out <= 16'hFFC8;    16'd48394: out <= 16'h016B;    16'd48395: out <= 16'h0158;
    16'd48396: out <= 16'h05E7;    16'd48397: out <= 16'h0077;    16'd48398: out <= 16'hFCA0;    16'd48399: out <= 16'hFD1A;
    16'd48400: out <= 16'hFEEE;    16'd48401: out <= 16'h0223;    16'd48402: out <= 16'h046C;    16'd48403: out <= 16'h05F1;
    16'd48404: out <= 16'h01C7;    16'd48405: out <= 16'h01CE;    16'd48406: out <= 16'hFF36;    16'd48407: out <= 16'hFD3F;
    16'd48408: out <= 16'h0104;    16'd48409: out <= 16'hFD7A;    16'd48410: out <= 16'hFC3D;    16'd48411: out <= 16'hFC89;
    16'd48412: out <= 16'h034D;    16'd48413: out <= 16'hFC85;    16'd48414: out <= 16'h01F3;    16'd48415: out <= 16'hFF2E;
    16'd48416: out <= 16'hFEA5;    16'd48417: out <= 16'hFE15;    16'd48418: out <= 16'h03AB;    16'd48419: out <= 16'hFC47;
    16'd48420: out <= 16'h00CF;    16'd48421: out <= 16'h0643;    16'd48422: out <= 16'hFB22;    16'd48423: out <= 16'h0452;
    16'd48424: out <= 16'h01CF;    16'd48425: out <= 16'h03C9;    16'd48426: out <= 16'h02D8;    16'd48427: out <= 16'h08AA;
    16'd48428: out <= 16'hFEF2;    16'd48429: out <= 16'h0616;    16'd48430: out <= 16'h0450;    16'd48431: out <= 16'h005C;
    16'd48432: out <= 16'h0260;    16'd48433: out <= 16'h07D4;    16'd48434: out <= 16'h00C8;    16'd48435: out <= 16'h0819;
    16'd48436: out <= 16'h0970;    16'd48437: out <= 16'h05FE;    16'd48438: out <= 16'h0301;    16'd48439: out <= 16'h02C9;
    16'd48440: out <= 16'h063B;    16'd48441: out <= 16'h019C;    16'd48442: out <= 16'hFFE4;    16'd48443: out <= 16'h032A;
    16'd48444: out <= 16'h043D;    16'd48445: out <= 16'h0171;    16'd48446: out <= 16'h01C0;    16'd48447: out <= 16'h04FF;
    16'd48448: out <= 16'h05D6;    16'd48449: out <= 16'hFCDA;    16'd48450: out <= 16'h0210;    16'd48451: out <= 16'hFFA8;
    16'd48452: out <= 16'h0434;    16'd48453: out <= 16'h0387;    16'd48454: out <= 16'h0BDE;    16'd48455: out <= 16'h014C;
    16'd48456: out <= 16'hFE16;    16'd48457: out <= 16'h07D2;    16'd48458: out <= 16'h0386;    16'd48459: out <= 16'h095F;
    16'd48460: out <= 16'h0995;    16'd48461: out <= 16'h0497;    16'd48462: out <= 16'hFB3E;    16'd48463: out <= 16'h0D84;
    16'd48464: out <= 16'h0061;    16'd48465: out <= 16'h006B;    16'd48466: out <= 16'h079B;    16'd48467: out <= 16'h00E6;
    16'd48468: out <= 16'h057E;    16'd48469: out <= 16'h0161;    16'd48470: out <= 16'h0A48;    16'd48471: out <= 16'h0153;
    16'd48472: out <= 16'h015C;    16'd48473: out <= 16'h0294;    16'd48474: out <= 16'h0481;    16'd48475: out <= 16'h01C6;
    16'd48476: out <= 16'h02CF;    16'd48477: out <= 16'h0742;    16'd48478: out <= 16'h0797;    16'd48479: out <= 16'h09C8;
    16'd48480: out <= 16'h03B8;    16'd48481: out <= 16'h0287;    16'd48482: out <= 16'hFB27;    16'd48483: out <= 16'h0CC0;
    16'd48484: out <= 16'h07EA;    16'd48485: out <= 16'hFFD4;    16'd48486: out <= 16'h069B;    16'd48487: out <= 16'h0AE3;
    16'd48488: out <= 16'h07C0;    16'd48489: out <= 16'h0563;    16'd48490: out <= 16'h0026;    16'd48491: out <= 16'hFF86;
    16'd48492: out <= 16'hFFF7;    16'd48493: out <= 16'hFF00;    16'd48494: out <= 16'hFB80;    16'd48495: out <= 16'h0C19;
    16'd48496: out <= 16'h067B;    16'd48497: out <= 16'hFDE9;    16'd48498: out <= 16'hFFC8;    16'd48499: out <= 16'h0572;
    16'd48500: out <= 16'hFD43;    16'd48501: out <= 16'hFF7D;    16'd48502: out <= 16'h0572;    16'd48503: out <= 16'h052F;
    16'd48504: out <= 16'h00B8;    16'd48505: out <= 16'h0147;    16'd48506: out <= 16'h043B;    16'd48507: out <= 16'h040A;
    16'd48508: out <= 16'h040B;    16'd48509: out <= 16'h04D3;    16'd48510: out <= 16'h0113;    16'd48511: out <= 16'h0139;
    16'd48512: out <= 16'h0825;    16'd48513: out <= 16'h051F;    16'd48514: out <= 16'h071A;    16'd48515: out <= 16'h0575;
    16'd48516: out <= 16'h04A6;    16'd48517: out <= 16'h0A02;    16'd48518: out <= 16'h020D;    16'd48519: out <= 16'h0820;
    16'd48520: out <= 16'h0383;    16'd48521: out <= 16'h0542;    16'd48522: out <= 16'h05C7;    16'd48523: out <= 16'h03C3;
    16'd48524: out <= 16'h0A5B;    16'd48525: out <= 16'hFA88;    16'd48526: out <= 16'h075A;    16'd48527: out <= 16'h00F4;
    16'd48528: out <= 16'h0601;    16'd48529: out <= 16'hFC8A;    16'd48530: out <= 16'h00E8;    16'd48531: out <= 16'h07C5;
    16'd48532: out <= 16'h05E2;    16'd48533: out <= 16'h08B9;    16'd48534: out <= 16'h08AE;    16'd48535: out <= 16'h04FB;
    16'd48536: out <= 16'hFF9E;    16'd48537: out <= 16'h04C3;    16'd48538: out <= 16'h02E8;    16'd48539: out <= 16'h0240;
    16'd48540: out <= 16'h017A;    16'd48541: out <= 16'h0206;    16'd48542: out <= 16'h02D8;    16'd48543: out <= 16'h037C;
    16'd48544: out <= 16'h0640;    16'd48545: out <= 16'h0AEB;    16'd48546: out <= 16'h0400;    16'd48547: out <= 16'h009A;
    16'd48548: out <= 16'hFFD6;    16'd48549: out <= 16'h0853;    16'd48550: out <= 16'h005C;    16'd48551: out <= 16'h0748;
    16'd48552: out <= 16'hFE14;    16'd48553: out <= 16'h0613;    16'd48554: out <= 16'h07AC;    16'd48555: out <= 16'h038A;
    16'd48556: out <= 16'h04CB;    16'd48557: out <= 16'h0907;    16'd48558: out <= 16'h0AA7;    16'd48559: out <= 16'h033F;
    16'd48560: out <= 16'h0B83;    16'd48561: out <= 16'h0947;    16'd48562: out <= 16'hFF4A;    16'd48563: out <= 16'h0186;
    16'd48564: out <= 16'hFF7F;    16'd48565: out <= 16'h063D;    16'd48566: out <= 16'h0742;    16'd48567: out <= 16'hFF2E;
    16'd48568: out <= 16'hFEE0;    16'd48569: out <= 16'h04CC;    16'd48570: out <= 16'h094E;    16'd48571: out <= 16'h055C;
    16'd48572: out <= 16'h010C;    16'd48573: out <= 16'h097C;    16'd48574: out <= 16'h0108;    16'd48575: out <= 16'h004E;
    16'd48576: out <= 16'h0A6A;    16'd48577: out <= 16'h0434;    16'd48578: out <= 16'h0330;    16'd48579: out <= 16'h06C9;
    16'd48580: out <= 16'h04DA;    16'd48581: out <= 16'h07CA;    16'd48582: out <= 16'hFB95;    16'd48583: out <= 16'h0484;
    16'd48584: out <= 16'h01AC;    16'd48585: out <= 16'hF6D1;    16'd48586: out <= 16'h01B0;    16'd48587: out <= 16'hFAFF;
    16'd48588: out <= 16'h0037;    16'd48589: out <= 16'hF8CA;    16'd48590: out <= 16'hFD82;    16'd48591: out <= 16'h009B;
    16'd48592: out <= 16'hFE07;    16'd48593: out <= 16'hFEE5;    16'd48594: out <= 16'hF868;    16'd48595: out <= 16'h04F9;
    16'd48596: out <= 16'hFCEC;    16'd48597: out <= 16'h0170;    16'd48598: out <= 16'hFB61;    16'd48599: out <= 16'h03DB;
    16'd48600: out <= 16'hFD16;    16'd48601: out <= 16'hFFA7;    16'd48602: out <= 16'h04B0;    16'd48603: out <= 16'h046F;
    16'd48604: out <= 16'h0423;    16'd48605: out <= 16'h05B6;    16'd48606: out <= 16'hFE17;    16'd48607: out <= 16'hFBB5;
    16'd48608: out <= 16'h00C3;    16'd48609: out <= 16'h02E1;    16'd48610: out <= 16'hFF6B;    16'd48611: out <= 16'hFE59;
    16'd48612: out <= 16'h02D5;    16'd48613: out <= 16'h0180;    16'd48614: out <= 16'hFEF0;    16'd48615: out <= 16'hFE8C;
    16'd48616: out <= 16'hFC38;    16'd48617: out <= 16'hFB99;    16'd48618: out <= 16'hFEB9;    16'd48619: out <= 16'h0250;
    16'd48620: out <= 16'hF7AE;    16'd48621: out <= 16'hFE22;    16'd48622: out <= 16'h0378;    16'd48623: out <= 16'h0282;
    16'd48624: out <= 16'hFFCD;    16'd48625: out <= 16'hFDA8;    16'd48626: out <= 16'hFFBE;    16'd48627: out <= 16'hFC68;
    16'd48628: out <= 16'h0954;    16'd48629: out <= 16'hFF9B;    16'd48630: out <= 16'hFF50;    16'd48631: out <= 16'hFC7E;
    16'd48632: out <= 16'hFC36;    16'd48633: out <= 16'h0341;    16'd48634: out <= 16'h018D;    16'd48635: out <= 16'hF7BC;
    16'd48636: out <= 16'h0938;    16'd48637: out <= 16'hFF4E;    16'd48638: out <= 16'hFEBC;    16'd48639: out <= 16'h02C3;
    16'd48640: out <= 16'hFED6;    16'd48641: out <= 16'hFD99;    16'd48642: out <= 16'hFDCB;    16'd48643: out <= 16'h009C;
    16'd48644: out <= 16'hFEA1;    16'd48645: out <= 16'hFDA4;    16'd48646: out <= 16'h00EE;    16'd48647: out <= 16'hFA16;
    16'd48648: out <= 16'h03BA;    16'd48649: out <= 16'h00D4;    16'd48650: out <= 16'h0220;    16'd48651: out <= 16'hFBFA;
    16'd48652: out <= 16'hFDAF;    16'd48653: out <= 16'h01D8;    16'd48654: out <= 16'h0066;    16'd48655: out <= 16'hFE3E;
    16'd48656: out <= 16'h016A;    16'd48657: out <= 16'h0372;    16'd48658: out <= 16'h0518;    16'd48659: out <= 16'h01C4;
    16'd48660: out <= 16'h0463;    16'd48661: out <= 16'h005E;    16'd48662: out <= 16'h02BF;    16'd48663: out <= 16'h0232;
    16'd48664: out <= 16'hF91A;    16'd48665: out <= 16'hFE83;    16'd48666: out <= 16'hFF64;    16'd48667: out <= 16'h0291;
    16'd48668: out <= 16'hFB1E;    16'd48669: out <= 16'hFB52;    16'd48670: out <= 16'hFEE2;    16'd48671: out <= 16'hFC17;
    16'd48672: out <= 16'h0297;    16'd48673: out <= 16'hFEDC;    16'd48674: out <= 16'h0006;    16'd48675: out <= 16'hFF23;
    16'd48676: out <= 16'hFC9C;    16'd48677: out <= 16'h01F0;    16'd48678: out <= 16'h0011;    16'd48679: out <= 16'h0471;
    16'd48680: out <= 16'h05B6;    16'd48681: out <= 16'h0307;    16'd48682: out <= 16'h00D4;    16'd48683: out <= 16'hFE50;
    16'd48684: out <= 16'h0AF8;    16'd48685: out <= 16'h03B1;    16'd48686: out <= 16'h0523;    16'd48687: out <= 16'h00C8;
    16'd48688: out <= 16'h01DC;    16'd48689: out <= 16'h056C;    16'd48690: out <= 16'h07C3;    16'd48691: out <= 16'h0254;
    16'd48692: out <= 16'h05F7;    16'd48693: out <= 16'h06DB;    16'd48694: out <= 16'h017F;    16'd48695: out <= 16'h01E3;
    16'd48696: out <= 16'h040B;    16'd48697: out <= 16'h079B;    16'd48698: out <= 16'h02A8;    16'd48699: out <= 16'h0618;
    16'd48700: out <= 16'h05DE;    16'd48701: out <= 16'h03CF;    16'd48702: out <= 16'h06BC;    16'd48703: out <= 16'h065E;
    16'd48704: out <= 16'h03FA;    16'd48705: out <= 16'h062A;    16'd48706: out <= 16'hFDF5;    16'd48707: out <= 16'h0B7E;
    16'd48708: out <= 16'hFEF4;    16'd48709: out <= 16'h057D;    16'd48710: out <= 16'h0092;    16'd48711: out <= 16'hFD15;
    16'd48712: out <= 16'h0062;    16'd48713: out <= 16'hFF74;    16'd48714: out <= 16'h015D;    16'd48715: out <= 16'h01DB;
    16'd48716: out <= 16'h0317;    16'd48717: out <= 16'h0585;    16'd48718: out <= 16'h09EB;    16'd48719: out <= 16'h0125;
    16'd48720: out <= 16'h0666;    16'd48721: out <= 16'h0B47;    16'd48722: out <= 16'h0B0E;    16'd48723: out <= 16'h0256;
    16'd48724: out <= 16'h0192;    16'd48725: out <= 16'h046A;    16'd48726: out <= 16'h0705;    16'd48727: out <= 16'hFFCF;
    16'd48728: out <= 16'h02DC;    16'd48729: out <= 16'h05B9;    16'd48730: out <= 16'hFF3D;    16'd48731: out <= 16'h004F;
    16'd48732: out <= 16'hFF5E;    16'd48733: out <= 16'h06B3;    16'd48734: out <= 16'h0938;    16'd48735: out <= 16'h0A8E;
    16'd48736: out <= 16'hFF0D;    16'd48737: out <= 16'h078C;    16'd48738: out <= 16'h0884;    16'd48739: out <= 16'h0167;
    16'd48740: out <= 16'h0144;    16'd48741: out <= 16'h062C;    16'd48742: out <= 16'h087C;    16'd48743: out <= 16'h03F4;
    16'd48744: out <= 16'h051F;    16'd48745: out <= 16'h068A;    16'd48746: out <= 16'h037E;    16'd48747: out <= 16'h0325;
    16'd48748: out <= 16'h095C;    16'd48749: out <= 16'h04FA;    16'd48750: out <= 16'h040A;    16'd48751: out <= 16'h01D5;
    16'd48752: out <= 16'h0349;    16'd48753: out <= 16'h04BC;    16'd48754: out <= 16'h075A;    16'd48755: out <= 16'h008A;
    16'd48756: out <= 16'h0A03;    16'd48757: out <= 16'h01F1;    16'd48758: out <= 16'h030A;    16'd48759: out <= 16'h02DB;
    16'd48760: out <= 16'h03B4;    16'd48761: out <= 16'h07FC;    16'd48762: out <= 16'h04DD;    16'd48763: out <= 16'h038E;
    16'd48764: out <= 16'h00B3;    16'd48765: out <= 16'hFFE3;    16'd48766: out <= 16'h07CD;    16'd48767: out <= 16'h07CB;
    16'd48768: out <= 16'h0572;    16'd48769: out <= 16'h03B0;    16'd48770: out <= 16'h03D0;    16'd48771: out <= 16'h041D;
    16'd48772: out <= 16'h0447;    16'd48773: out <= 16'h06B9;    16'd48774: out <= 16'h0B7E;    16'd48775: out <= 16'h06D2;
    16'd48776: out <= 16'h0518;    16'd48777: out <= 16'h02FA;    16'd48778: out <= 16'h007B;    16'd48779: out <= 16'hFE02;
    16'd48780: out <= 16'h04CC;    16'd48781: out <= 16'h021B;    16'd48782: out <= 16'h05CF;    16'd48783: out <= 16'h017F;
    16'd48784: out <= 16'h015E;    16'd48785: out <= 16'h052C;    16'd48786: out <= 16'h003C;    16'd48787: out <= 16'h006B;
    16'd48788: out <= 16'h0768;    16'd48789: out <= 16'h045C;    16'd48790: out <= 16'h0D99;    16'd48791: out <= 16'h0175;
    16'd48792: out <= 16'h05E9;    16'd48793: out <= 16'h0A01;    16'd48794: out <= 16'h0197;    16'd48795: out <= 16'h0D4C;
    16'd48796: out <= 16'h07A5;    16'd48797: out <= 16'h0209;    16'd48798: out <= 16'h06EC;    16'd48799: out <= 16'h0966;
    16'd48800: out <= 16'h0E52;    16'd48801: out <= 16'h0265;    16'd48802: out <= 16'h0837;    16'd48803: out <= 16'hFF56;
    16'd48804: out <= 16'h05BC;    16'd48805: out <= 16'h0C6E;    16'd48806: out <= 16'h0327;    16'd48807: out <= 16'h0012;
    16'd48808: out <= 16'h0EFD;    16'd48809: out <= 16'h04A1;    16'd48810: out <= 16'h0712;    16'd48811: out <= 16'h07A4;
    16'd48812: out <= 16'hFD40;    16'd48813: out <= 16'h05AD;    16'd48814: out <= 16'hFDBE;    16'd48815: out <= 16'h0272;
    16'd48816: out <= 16'h09DC;    16'd48817: out <= 16'h0BD8;    16'd48818: out <= 16'h0900;    16'd48819: out <= 16'hFB26;
    16'd48820: out <= 16'h0451;    16'd48821: out <= 16'h0546;    16'd48822: out <= 16'h044A;    16'd48823: out <= 16'h028B;
    16'd48824: out <= 16'h0358;    16'd48825: out <= 16'h051E;    16'd48826: out <= 16'h03EC;    16'd48827: out <= 16'h0844;
    16'd48828: out <= 16'h0255;    16'd48829: out <= 16'h00AA;    16'd48830: out <= 16'hFE3D;    16'd48831: out <= 16'h00CB;
    16'd48832: out <= 16'h026A;    16'd48833: out <= 16'h080D;    16'd48834: out <= 16'h0343;    16'd48835: out <= 16'h0112;
    16'd48836: out <= 16'h04B5;    16'd48837: out <= 16'h0366;    16'd48838: out <= 16'hFE4C;    16'd48839: out <= 16'hFFF1;
    16'd48840: out <= 16'h03C0;    16'd48841: out <= 16'h0460;    16'd48842: out <= 16'hF668;    16'd48843: out <= 16'h09AB;
    16'd48844: out <= 16'hFF61;    16'd48845: out <= 16'h02D9;    16'd48846: out <= 16'hF97D;    16'd48847: out <= 16'h04D5;
    16'd48848: out <= 16'h0136;    16'd48849: out <= 16'h0200;    16'd48850: out <= 16'h00CA;    16'd48851: out <= 16'hFDF8;
    16'd48852: out <= 16'h06A9;    16'd48853: out <= 16'hFF12;    16'd48854: out <= 16'hFED8;    16'd48855: out <= 16'hFD2D;
    16'd48856: out <= 16'hFF2D;    16'd48857: out <= 16'h033C;    16'd48858: out <= 16'h004F;    16'd48859: out <= 16'hFE6E;
    16'd48860: out <= 16'hFF6A;    16'd48861: out <= 16'h00E0;    16'd48862: out <= 16'hFDE1;    16'd48863: out <= 16'h020E;
    16'd48864: out <= 16'h000B;    16'd48865: out <= 16'hF95D;    16'd48866: out <= 16'hFFEF;    16'd48867: out <= 16'hFD7B;
    16'd48868: out <= 16'hFE9D;    16'd48869: out <= 16'h036F;    16'd48870: out <= 16'h0574;    16'd48871: out <= 16'hF930;
    16'd48872: out <= 16'h04DE;    16'd48873: out <= 16'h04CC;    16'd48874: out <= 16'hFC37;    16'd48875: out <= 16'h0524;
    16'd48876: out <= 16'hF570;    16'd48877: out <= 16'h0266;    16'd48878: out <= 16'hFCF5;    16'd48879: out <= 16'hFDD0;
    16'd48880: out <= 16'hFDAB;    16'd48881: out <= 16'h0572;    16'd48882: out <= 16'hFA5C;    16'd48883: out <= 16'hFCAA;
    16'd48884: out <= 16'h032B;    16'd48885: out <= 16'hFFC0;    16'd48886: out <= 16'h00B1;    16'd48887: out <= 16'h03C7;
    16'd48888: out <= 16'h014A;    16'd48889: out <= 16'hF99E;    16'd48890: out <= 16'hFD58;    16'd48891: out <= 16'hF96A;
    16'd48892: out <= 16'hFF03;    16'd48893: out <= 16'hFF97;    16'd48894: out <= 16'h0557;    16'd48895: out <= 16'hFE9D;
    16'd48896: out <= 16'h0159;    16'd48897: out <= 16'hFB77;    16'd48898: out <= 16'hF7EC;    16'd48899: out <= 16'h0246;
    16'd48900: out <= 16'hF995;    16'd48901: out <= 16'h04E3;    16'd48902: out <= 16'hFB91;    16'd48903: out <= 16'h0062;
    16'd48904: out <= 16'h0454;    16'd48905: out <= 16'h0154;    16'd48906: out <= 16'h0357;    16'd48907: out <= 16'hFF53;
    16'd48908: out <= 16'hFE79;    16'd48909: out <= 16'hFB4B;    16'd48910: out <= 16'h00A5;    16'd48911: out <= 16'h0445;
    16'd48912: out <= 16'hFCCE;    16'd48913: out <= 16'h033A;    16'd48914: out <= 16'hFD7A;    16'd48915: out <= 16'h0156;
    16'd48916: out <= 16'hFC8A;    16'd48917: out <= 16'h0239;    16'd48918: out <= 16'hFEAC;    16'd48919: out <= 16'h00F1;
    16'd48920: out <= 16'hFB29;    16'd48921: out <= 16'h0052;    16'd48922: out <= 16'h012F;    16'd48923: out <= 16'hFC1D;
    16'd48924: out <= 16'hFFD7;    16'd48925: out <= 16'h0155;    16'd48926: out <= 16'hFF10;    16'd48927: out <= 16'hF9DA;
    16'd48928: out <= 16'h0577;    16'd48929: out <= 16'hFF13;    16'd48930: out <= 16'h0034;    16'd48931: out <= 16'h016A;
    16'd48932: out <= 16'hFA2E;    16'd48933: out <= 16'h0250;    16'd48934: out <= 16'hFD96;    16'd48935: out <= 16'hF90B;
    16'd48936: out <= 16'hFDAD;    16'd48937: out <= 16'h0574;    16'd48938: out <= 16'h0811;    16'd48939: out <= 16'h0AA4;
    16'd48940: out <= 16'h0189;    16'd48941: out <= 16'h04DF;    16'd48942: out <= 16'h05AF;    16'd48943: out <= 16'hFBE8;
    16'd48944: out <= 16'h081F;    16'd48945: out <= 16'h0B3C;    16'd48946: out <= 16'hFE21;    16'd48947: out <= 16'h04B8;
    16'd48948: out <= 16'hFD2C;    16'd48949: out <= 16'h02ED;    16'd48950: out <= 16'hFF43;    16'd48951: out <= 16'h03C6;
    16'd48952: out <= 16'h02B4;    16'd48953: out <= 16'h0623;    16'd48954: out <= 16'h0109;    16'd48955: out <= 16'h0848;
    16'd48956: out <= 16'h01A3;    16'd48957: out <= 16'h069C;    16'd48958: out <= 16'h0114;    16'd48959: out <= 16'h0320;
    16'd48960: out <= 16'h0578;    16'd48961: out <= 16'h0858;    16'd48962: out <= 16'h0531;    16'd48963: out <= 16'h0298;
    16'd48964: out <= 16'h017B;    16'd48965: out <= 16'h02F7;    16'd48966: out <= 16'h05BA;    16'd48967: out <= 16'h0732;
    16'd48968: out <= 16'h05EF;    16'd48969: out <= 16'h018A;    16'd48970: out <= 16'h0223;    16'd48971: out <= 16'h0373;
    16'd48972: out <= 16'h014F;    16'd48973: out <= 16'h0459;    16'd48974: out <= 16'h02E8;    16'd48975: out <= 16'h0513;
    16'd48976: out <= 16'h07C3;    16'd48977: out <= 16'h0A93;    16'd48978: out <= 16'hFE24;    16'd48979: out <= 16'h07C2;
    16'd48980: out <= 16'h0484;    16'd48981: out <= 16'h0455;    16'd48982: out <= 16'h042D;    16'd48983: out <= 16'h0521;
    16'd48984: out <= 16'h053B;    16'd48985: out <= 16'h07A3;    16'd48986: out <= 16'h05A1;    16'd48987: out <= 16'h0533;
    16'd48988: out <= 16'hFCD2;    16'd48989: out <= 16'h08AB;    16'd48990: out <= 16'hFAA7;    16'd48991: out <= 16'h0265;
    16'd48992: out <= 16'h0C13;    16'd48993: out <= 16'h0225;    16'd48994: out <= 16'h02D6;    16'd48995: out <= 16'h0534;
    16'd48996: out <= 16'h04F0;    16'd48997: out <= 16'h0625;    16'd48998: out <= 16'h0647;    16'd48999: out <= 16'h035B;
    16'd49000: out <= 16'h07F5;    16'd49001: out <= 16'h03F6;    16'd49002: out <= 16'h03BD;    16'd49003: out <= 16'h084D;
    16'd49004: out <= 16'h07AD;    16'd49005: out <= 16'hFE99;    16'd49006: out <= 16'hFE54;    16'd49007: out <= 16'h05B5;
    16'd49008: out <= 16'hFF08;    16'd49009: out <= 16'h0389;    16'd49010: out <= 16'h008E;    16'd49011: out <= 16'h06D9;
    16'd49012: out <= 16'h06F4;    16'd49013: out <= 16'hFD35;    16'd49014: out <= 16'hFF59;    16'd49015: out <= 16'h076F;
    16'd49016: out <= 16'h05A6;    16'd49017: out <= 16'h01F9;    16'd49018: out <= 16'h0235;    16'd49019: out <= 16'h0353;
    16'd49020: out <= 16'h0000;    16'd49021: out <= 16'h0B71;    16'd49022: out <= 16'h08AD;    16'd49023: out <= 16'h0625;
    16'd49024: out <= 16'h01D1;    16'd49025: out <= 16'hFD6E;    16'd49026: out <= 16'h042B;    16'd49027: out <= 16'h05A3;
    16'd49028: out <= 16'h07C8;    16'd49029: out <= 16'h0536;    16'd49030: out <= 16'h038C;    16'd49031: out <= 16'h0201;
    16'd49032: out <= 16'h055A;    16'd49033: out <= 16'h027D;    16'd49034: out <= 16'h0B03;    16'd49035: out <= 16'hFF0C;
    16'd49036: out <= 16'hFFBB;    16'd49037: out <= 16'h0208;    16'd49038: out <= 16'h0893;    16'd49039: out <= 16'hFD27;
    16'd49040: out <= 16'h04E3;    16'd49041: out <= 16'hFF72;    16'd49042: out <= 16'h0039;    16'd49043: out <= 16'h08B7;
    16'd49044: out <= 16'h03E5;    16'd49045: out <= 16'h07AD;    16'd49046: out <= 16'h061D;    16'd49047: out <= 16'h06CA;
    16'd49048: out <= 16'h0191;    16'd49049: out <= 16'h0D60;    16'd49050: out <= 16'h0BA8;    16'd49051: out <= 16'h07A8;
    16'd49052: out <= 16'h03CD;    16'd49053: out <= 16'hFF3D;    16'd49054: out <= 16'h079E;    16'd49055: out <= 16'hFF6E;
    16'd49056: out <= 16'hFEC4;    16'd49057: out <= 16'h045B;    16'd49058: out <= 16'h0433;    16'd49059: out <= 16'h0065;
    16'd49060: out <= 16'h065A;    16'd49061: out <= 16'h00A0;    16'd49062: out <= 16'h095F;    16'd49063: out <= 16'h000E;
    16'd49064: out <= 16'h02D5;    16'd49065: out <= 16'h0700;    16'd49066: out <= 16'h02BA;    16'd49067: out <= 16'h03FF;
    16'd49068: out <= 16'h0696;    16'd49069: out <= 16'hFA8F;    16'd49070: out <= 16'h0074;    16'd49071: out <= 16'h03C7;
    16'd49072: out <= 16'h04EF;    16'd49073: out <= 16'h0CC2;    16'd49074: out <= 16'h0AF4;    16'd49075: out <= 16'h0804;
    16'd49076: out <= 16'h01FF;    16'd49077: out <= 16'h0523;    16'd49078: out <= 16'hFFFF;    16'd49079: out <= 16'h0018;
    16'd49080: out <= 16'h03C4;    16'd49081: out <= 16'h0336;    16'd49082: out <= 16'h03FF;    16'd49083: out <= 16'h07E5;
    16'd49084: out <= 16'h00D4;    16'd49085: out <= 16'h08E9;    16'd49086: out <= 16'h0474;    16'd49087: out <= 16'h0478;
    16'd49088: out <= 16'h05A7;    16'd49089: out <= 16'h080A;    16'd49090: out <= 16'h0780;    16'd49091: out <= 16'hFFBF;
    16'd49092: out <= 16'h06DF;    16'd49093: out <= 16'hFD08;    16'd49094: out <= 16'h00E9;    16'd49095: out <= 16'hFEA1;
    16'd49096: out <= 16'hFBE9;    16'd49097: out <= 16'h0248;    16'd49098: out <= 16'hFE82;    16'd49099: out <= 16'hFD02;
    16'd49100: out <= 16'hFE37;    16'd49101: out <= 16'hFD07;    16'd49102: out <= 16'hF711;    16'd49103: out <= 16'hFC0F;
    16'd49104: out <= 16'hFDA1;    16'd49105: out <= 16'hFEE1;    16'd49106: out <= 16'h01D5;    16'd49107: out <= 16'h041C;
    16'd49108: out <= 16'h0041;    16'd49109: out <= 16'hFD60;    16'd49110: out <= 16'hFDE7;    16'd49111: out <= 16'h0123;
    16'd49112: out <= 16'hFB5E;    16'd49113: out <= 16'hF91F;    16'd49114: out <= 16'h0148;    16'd49115: out <= 16'hFCC6;
    16'd49116: out <= 16'hFF6A;    16'd49117: out <= 16'h048E;    16'd49118: out <= 16'h04D4;    16'd49119: out <= 16'hFED3;
    16'd49120: out <= 16'h0430;    16'd49121: out <= 16'h01D3;    16'd49122: out <= 16'hFC4B;    16'd49123: out <= 16'hFE3B;
    16'd49124: out <= 16'h011B;    16'd49125: out <= 16'h00B5;    16'd49126: out <= 16'hF7EC;    16'd49127: out <= 16'h05D5;
    16'd49128: out <= 16'h011B;    16'd49129: out <= 16'h02E5;    16'd49130: out <= 16'h0384;    16'd49131: out <= 16'hFAEB;
    16'd49132: out <= 16'hF7FC;    16'd49133: out <= 16'h02D7;    16'd49134: out <= 16'h021B;    16'd49135: out <= 16'hFDBA;
    16'd49136: out <= 16'h000B;    16'd49137: out <= 16'hF8A8;    16'd49138: out <= 16'h046D;    16'd49139: out <= 16'h01D7;
    16'd49140: out <= 16'h01B3;    16'd49141: out <= 16'h01F1;    16'd49142: out <= 16'hFC10;    16'd49143: out <= 16'hFD16;
    16'd49144: out <= 16'hFDC9;    16'd49145: out <= 16'h0290;    16'd49146: out <= 16'hFE84;    16'd49147: out <= 16'h02C2;
    16'd49148: out <= 16'hFE2D;    16'd49149: out <= 16'hF87A;    16'd49150: out <= 16'hF9EE;    16'd49151: out <= 16'h0464;
    16'd49152: out <= 16'h00EE;    16'd49153: out <= 16'h01D8;    16'd49154: out <= 16'h02BD;    16'd49155: out <= 16'h0003;
    16'd49156: out <= 16'h00C8;    16'd49157: out <= 16'h035F;    16'd49158: out <= 16'h00DE;    16'd49159: out <= 16'hFD86;
    16'd49160: out <= 16'hFE1D;    16'd49161: out <= 16'hFDCE;    16'd49162: out <= 16'hFFA2;    16'd49163: out <= 16'h0323;
    16'd49164: out <= 16'h0354;    16'd49165: out <= 16'h08B4;    16'd49166: out <= 16'hFF68;    16'd49167: out <= 16'hFEAC;
    16'd49168: out <= 16'h0418;    16'd49169: out <= 16'hFABB;    16'd49170: out <= 16'hFE26;    16'd49171: out <= 16'hFACF;
    16'd49172: out <= 16'hFBC3;    16'd49173: out <= 16'hFFCF;    16'd49174: out <= 16'h02F1;    16'd49175: out <= 16'hFAF6;
    16'd49176: out <= 16'hFA4E;    16'd49177: out <= 16'h028C;    16'd49178: out <= 16'h03BE;    16'd49179: out <= 16'h05D3;
    16'd49180: out <= 16'h01BB;    16'd49181: out <= 16'h08DD;    16'd49182: out <= 16'hFB4C;    16'd49183: out <= 16'h038D;
    16'd49184: out <= 16'h0496;    16'd49185: out <= 16'h05F7;    16'd49186: out <= 16'h009E;    16'd49187: out <= 16'h040A;
    16'd49188: out <= 16'h018B;    16'd49189: out <= 16'hF906;    16'd49190: out <= 16'h02B7;    16'd49191: out <= 16'h04E6;
    16'd49192: out <= 16'h01CA;    16'd49193: out <= 16'h0934;    16'd49194: out <= 16'h0580;    16'd49195: out <= 16'h033C;
    16'd49196: out <= 16'h0821;    16'd49197: out <= 16'h0307;    16'd49198: out <= 16'h0508;    16'd49199: out <= 16'h0A36;
    16'd49200: out <= 16'h00B5;    16'd49201: out <= 16'h050D;    16'd49202: out <= 16'h006C;    16'd49203: out <= 16'hFA7E;
    16'd49204: out <= 16'h0150;    16'd49205: out <= 16'h08D2;    16'd49206: out <= 16'h028B;    16'd49207: out <= 16'h05D7;
    16'd49208: out <= 16'h013D;    16'd49209: out <= 16'h0487;    16'd49210: out <= 16'hFA1A;    16'd49211: out <= 16'h08DE;
    16'd49212: out <= 16'h02ED;    16'd49213: out <= 16'h02DE;    16'd49214: out <= 16'h036E;    16'd49215: out <= 16'h00DE;
    16'd49216: out <= 16'h0B0B;    16'd49217: out <= 16'h0087;    16'd49218: out <= 16'h0996;    16'd49219: out <= 16'h0352;
    16'd49220: out <= 16'h00DA;    16'd49221: out <= 16'h0873;    16'd49222: out <= 16'h0326;    16'd49223: out <= 16'hFE9A;
    16'd49224: out <= 16'h01B5;    16'd49225: out <= 16'h048B;    16'd49226: out <= 16'h0411;    16'd49227: out <= 16'h0AA6;
    16'd49228: out <= 16'h03F0;    16'd49229: out <= 16'h00F2;    16'd49230: out <= 16'h06B9;    16'd49231: out <= 16'h0628;
    16'd49232: out <= 16'h0A1B;    16'd49233: out <= 16'hFE26;    16'd49234: out <= 16'h06FB;    16'd49235: out <= 16'h0188;
    16'd49236: out <= 16'h0457;    16'd49237: out <= 16'h04D2;    16'd49238: out <= 16'h0751;    16'd49239: out <= 16'hFF90;
    16'd49240: out <= 16'hFEE4;    16'd49241: out <= 16'hFCD4;    16'd49242: out <= 16'h0738;    16'd49243: out <= 16'h07F5;
    16'd49244: out <= 16'h034C;    16'd49245: out <= 16'h0365;    16'd49246: out <= 16'h0351;    16'd49247: out <= 16'h068C;
    16'd49248: out <= 16'h06CB;    16'd49249: out <= 16'h0664;    16'd49250: out <= 16'h0886;    16'd49251: out <= 16'h0BDF;
    16'd49252: out <= 16'h0A24;    16'd49253: out <= 16'h01E8;    16'd49254: out <= 16'h0486;    16'd49255: out <= 16'h01C7;
    16'd49256: out <= 16'h02E9;    16'd49257: out <= 16'h0270;    16'd49258: out <= 16'h018C;    16'd49259: out <= 16'h04EC;
    16'd49260: out <= 16'h0826;    16'd49261: out <= 16'h00A5;    16'd49262: out <= 16'h073B;    16'd49263: out <= 16'h05C1;
    16'd49264: out <= 16'h028C;    16'd49265: out <= 16'h06D1;    16'd49266: out <= 16'h092F;    16'd49267: out <= 16'h0384;
    16'd49268: out <= 16'h0361;    16'd49269: out <= 16'h0486;    16'd49270: out <= 16'h0859;    16'd49271: out <= 16'h059F;
    16'd49272: out <= 16'hFFCA;    16'd49273: out <= 16'h017A;    16'd49274: out <= 16'h0656;    16'd49275: out <= 16'h02B0;
    16'd49276: out <= 16'h0395;    16'd49277: out <= 16'h018E;    16'd49278: out <= 16'hFD68;    16'd49279: out <= 16'h0664;
    16'd49280: out <= 16'h0755;    16'd49281: out <= 16'h036F;    16'd49282: out <= 16'h029B;    16'd49283: out <= 16'hFD28;
    16'd49284: out <= 16'h0656;    16'd49285: out <= 16'h06A0;    16'd49286: out <= 16'h0580;    16'd49287: out <= 16'h0005;
    16'd49288: out <= 16'hFECD;    16'd49289: out <= 16'h0420;    16'd49290: out <= 16'h026A;    16'd49291: out <= 16'hFEA4;
    16'd49292: out <= 16'hFBD2;    16'd49293: out <= 16'h00F8;    16'd49294: out <= 16'hFB97;    16'd49295: out <= 16'h0776;
    16'd49296: out <= 16'h05AC;    16'd49297: out <= 16'h01F5;    16'd49298: out <= 16'h057D;    16'd49299: out <= 16'h023F;
    16'd49300: out <= 16'hFF4C;    16'd49301: out <= 16'h055E;    16'd49302: out <= 16'h0600;    16'd49303: out <= 16'h027C;
    16'd49304: out <= 16'h005C;    16'd49305: out <= 16'h0591;    16'd49306: out <= 16'h09FC;    16'd49307: out <= 16'hFE1A;
    16'd49308: out <= 16'h0E53;    16'd49309: out <= 16'h073E;    16'd49310: out <= 16'h0382;    16'd49311: out <= 16'h0244;
    16'd49312: out <= 16'h06D6;    16'd49313: out <= 16'h0B2F;    16'd49314: out <= 16'h053F;    16'd49315: out <= 16'h05E4;
    16'd49316: out <= 16'h03F6;    16'd49317: out <= 16'h0326;    16'd49318: out <= 16'h07FF;    16'd49319: out <= 16'hFB0D;
    16'd49320: out <= 16'hFB24;    16'd49321: out <= 16'h1095;    16'd49322: out <= 16'h02DE;    16'd49323: out <= 16'h05A8;
    16'd49324: out <= 16'h0418;    16'd49325: out <= 16'h054E;    16'd49326: out <= 16'h0094;    16'd49327: out <= 16'hFFCA;
    16'd49328: out <= 16'h03F9;    16'd49329: out <= 16'h06A9;    16'd49330: out <= 16'h051D;    16'd49331: out <= 16'h023A;
    16'd49332: out <= 16'h06E3;    16'd49333: out <= 16'h086B;    16'd49334: out <= 16'hF89E;    16'd49335: out <= 16'h077D;
    16'd49336: out <= 16'h04D6;    16'd49337: out <= 16'hFAD7;    16'd49338: out <= 16'h029E;    16'd49339: out <= 16'h07E5;
    16'd49340: out <= 16'h015A;    16'd49341: out <= 16'h02B6;    16'd49342: out <= 16'h0197;    16'd49343: out <= 16'h047D;
    16'd49344: out <= 16'h0007;    16'd49345: out <= 16'h0256;    16'd49346: out <= 16'h0853;    16'd49347: out <= 16'h0144;
    16'd49348: out <= 16'hFE8F;    16'd49349: out <= 16'h0334;    16'd49350: out <= 16'hFEC5;    16'd49351: out <= 16'hFD39;
    16'd49352: out <= 16'hF8F5;    16'd49353: out <= 16'h070E;    16'd49354: out <= 16'h0368;    16'd49355: out <= 16'h0204;
    16'd49356: out <= 16'h0405;    16'd49357: out <= 16'h0045;    16'd49358: out <= 16'hFC75;    16'd49359: out <= 16'hFE8C;
    16'd49360: out <= 16'h025B;    16'd49361: out <= 16'hFE14;    16'd49362: out <= 16'h0039;    16'd49363: out <= 16'hFC31;
    16'd49364: out <= 16'hFD43;    16'd49365: out <= 16'h01D9;    16'd49366: out <= 16'hFE0E;    16'd49367: out <= 16'hFF2E;
    16'd49368: out <= 16'hFD69;    16'd49369: out <= 16'h051C;    16'd49370: out <= 16'hF7DD;    16'd49371: out <= 16'h0623;
    16'd49372: out <= 16'h01F0;    16'd49373: out <= 16'hFD71;    16'd49374: out <= 16'h01B3;    16'd49375: out <= 16'h049E;
    16'd49376: out <= 16'h0170;    16'd49377: out <= 16'hFD4B;    16'd49378: out <= 16'h019A;    16'd49379: out <= 16'hFD35;
    16'd49380: out <= 16'hFBAD;    16'd49381: out <= 16'h0702;    16'd49382: out <= 16'hFC72;    16'd49383: out <= 16'hFAF9;
    16'd49384: out <= 16'hFDC1;    16'd49385: out <= 16'h0218;    16'd49386: out <= 16'hFBA3;    16'd49387: out <= 16'h0135;
    16'd49388: out <= 16'h05C1;    16'd49389: out <= 16'h02C7;    16'd49390: out <= 16'hFD1A;    16'd49391: out <= 16'h033D;
    16'd49392: out <= 16'h0209;    16'd49393: out <= 16'h018D;    16'd49394: out <= 16'hFF58;    16'd49395: out <= 16'hF847;
    16'd49396: out <= 16'hFF54;    16'd49397: out <= 16'hFF2D;    16'd49398: out <= 16'hFE83;    16'd49399: out <= 16'hFF4D;
    16'd49400: out <= 16'h03BD;    16'd49401: out <= 16'h0BC6;    16'd49402: out <= 16'hFBC4;    16'd49403: out <= 16'hF941;
    16'd49404: out <= 16'h058B;    16'd49405: out <= 16'hFB14;    16'd49406: out <= 16'hFD7A;    16'd49407: out <= 16'h03F4;
    16'd49408: out <= 16'h035C;    16'd49409: out <= 16'h000A;    16'd49410: out <= 16'h03AC;    16'd49411: out <= 16'hFA78;
    16'd49412: out <= 16'h02BF;    16'd49413: out <= 16'h0027;    16'd49414: out <= 16'hFEAD;    16'd49415: out <= 16'h07D0;
    16'd49416: out <= 16'hFCA5;    16'd49417: out <= 16'h04DC;    16'd49418: out <= 16'hFFDE;    16'd49419: out <= 16'hFA80;
    16'd49420: out <= 16'hFDA8;    16'd49421: out <= 16'hFB60;    16'd49422: out <= 16'hFD4E;    16'd49423: out <= 16'h01F3;
    16'd49424: out <= 16'hFDCC;    16'd49425: out <= 16'hFD42;    16'd49426: out <= 16'h0497;    16'd49427: out <= 16'hFB3D;
    16'd49428: out <= 16'hFE19;    16'd49429: out <= 16'h0326;    16'd49430: out <= 16'hFADE;    16'd49431: out <= 16'h0372;
    16'd49432: out <= 16'hFB34;    16'd49433: out <= 16'h02C3;    16'd49434: out <= 16'hFC7C;    16'd49435: out <= 16'h06C9;
    16'd49436: out <= 16'hFF95;    16'd49437: out <= 16'hFA8E;    16'd49438: out <= 16'h051F;    16'd49439: out <= 16'hFEEF;
    16'd49440: out <= 16'h044F;    16'd49441: out <= 16'h03FA;    16'd49442: out <= 16'hFD5E;    16'd49443: out <= 16'hF9E5;
    16'd49444: out <= 16'hFEB7;    16'd49445: out <= 16'h05B7;    16'd49446: out <= 16'h006A;    16'd49447: out <= 16'hFD89;
    16'd49448: out <= 16'hFC98;    16'd49449: out <= 16'h0310;    16'd49450: out <= 16'hFDE8;    16'd49451: out <= 16'h0380;
    16'd49452: out <= 16'hFD44;    16'd49453: out <= 16'hFA74;    16'd49454: out <= 16'h06A2;    16'd49455: out <= 16'hFF9F;
    16'd49456: out <= 16'h03FE;    16'd49457: out <= 16'h02A8;    16'd49458: out <= 16'h07C0;    16'd49459: out <= 16'h0381;
    16'd49460: out <= 16'h032D;    16'd49461: out <= 16'h0570;    16'd49462: out <= 16'h0A6C;    16'd49463: out <= 16'h00C2;
    16'd49464: out <= 16'hFE0D;    16'd49465: out <= 16'h059A;    16'd49466: out <= 16'h0487;    16'd49467: out <= 16'h039A;
    16'd49468: out <= 16'h07D5;    16'd49469: out <= 16'h05A9;    16'd49470: out <= 16'h03AF;    16'd49471: out <= 16'h083F;
    16'd49472: out <= 16'hFE48;    16'd49473: out <= 16'h07FC;    16'd49474: out <= 16'h022F;    16'd49475: out <= 16'h05A3;
    16'd49476: out <= 16'h071C;    16'd49477: out <= 16'h0440;    16'd49478: out <= 16'h031A;    16'd49479: out <= 16'h0207;
    16'd49480: out <= 16'hFEE0;    16'd49481: out <= 16'h0034;    16'd49482: out <= 16'h03A6;    16'd49483: out <= 16'h04EE;
    16'd49484: out <= 16'h034E;    16'd49485: out <= 16'h02A8;    16'd49486: out <= 16'h050F;    16'd49487: out <= 16'h04D5;
    16'd49488: out <= 16'h08F8;    16'd49489: out <= 16'hFD30;    16'd49490: out <= 16'h09EA;    16'd49491: out <= 16'h041A;
    16'd49492: out <= 16'h04FD;    16'd49493: out <= 16'h0610;    16'd49494: out <= 16'h0727;    16'd49495: out <= 16'h059B;
    16'd49496: out <= 16'h0424;    16'd49497: out <= 16'h0B0F;    16'd49498: out <= 16'h04F7;    16'd49499: out <= 16'h0071;
    16'd49500: out <= 16'h0864;    16'd49501: out <= 16'h01F7;    16'd49502: out <= 16'h047E;    16'd49503: out <= 16'h0354;
    16'd49504: out <= 16'h0576;    16'd49505: out <= 16'h0887;    16'd49506: out <= 16'hFE95;    16'd49507: out <= 16'h0190;
    16'd49508: out <= 16'h0277;    16'd49509: out <= 16'h0321;    16'd49510: out <= 16'h0394;    16'd49511: out <= 16'h0380;
    16'd49512: out <= 16'h0514;    16'd49513: out <= 16'h029C;    16'd49514: out <= 16'h01FA;    16'd49515: out <= 16'hFD5E;
    16'd49516: out <= 16'h0271;    16'd49517: out <= 16'h00E2;    16'd49518: out <= 16'h0165;    16'd49519: out <= 16'h00AC;
    16'd49520: out <= 16'h07D1;    16'd49521: out <= 16'h062A;    16'd49522: out <= 16'h060D;    16'd49523: out <= 16'h0A68;
    16'd49524: out <= 16'hFEFB;    16'd49525: out <= 16'h05E5;    16'd49526: out <= 16'h017F;    16'd49527: out <= 16'h0243;
    16'd49528: out <= 16'hFE6D;    16'd49529: out <= 16'h06F2;    16'd49530: out <= 16'h007C;    16'd49531: out <= 16'h03EC;
    16'd49532: out <= 16'h03CE;    16'd49533: out <= 16'h06F7;    16'd49534: out <= 16'h0975;    16'd49535: out <= 16'hFE42;
    16'd49536: out <= 16'h01AD;    16'd49537: out <= 16'h004C;    16'd49538: out <= 16'hFF57;    16'd49539: out <= 16'h045E;
    16'd49540: out <= 16'hFD9B;    16'd49541: out <= 16'h0229;    16'd49542: out <= 16'h0522;    16'd49543: out <= 16'h03EB;
    16'd49544: out <= 16'h02CC;    16'd49545: out <= 16'h0477;    16'd49546: out <= 16'h02BF;    16'd49547: out <= 16'h03D2;
    16'd49548: out <= 16'h049A;    16'd49549: out <= 16'h048F;    16'd49550: out <= 16'h02A0;    16'd49551: out <= 16'h04E8;
    16'd49552: out <= 16'h0245;    16'd49553: out <= 16'h01ED;    16'd49554: out <= 16'h0479;    16'd49555: out <= 16'h05CF;
    16'd49556: out <= 16'h0B09;    16'd49557: out <= 16'h0153;    16'd49558: out <= 16'h078D;    16'd49559: out <= 16'h018A;
    16'd49560: out <= 16'h040F;    16'd49561: out <= 16'h0370;    16'd49562: out <= 16'h0385;    16'd49563: out <= 16'hFF3B;
    16'd49564: out <= 16'h00AE;    16'd49565: out <= 16'h067C;    16'd49566: out <= 16'h0130;    16'd49567: out <= 16'h020E;
    16'd49568: out <= 16'h05AF;    16'd49569: out <= 16'h0129;    16'd49570: out <= 16'h05A0;    16'd49571: out <= 16'h0502;
    16'd49572: out <= 16'h0504;    16'd49573: out <= 16'h02B9;    16'd49574: out <= 16'hFEA3;    16'd49575: out <= 16'h0618;
    16'd49576: out <= 16'h03CB;    16'd49577: out <= 16'h018B;    16'd49578: out <= 16'h02FF;    16'd49579: out <= 16'hFE6C;
    16'd49580: out <= 16'hFFAB;    16'd49581: out <= 16'h01DB;    16'd49582: out <= 16'h03A0;    16'd49583: out <= 16'h058B;
    16'd49584: out <= 16'h063C;    16'd49585: out <= 16'h0352;    16'd49586: out <= 16'h055A;    16'd49587: out <= 16'h052E;
    16'd49588: out <= 16'h076C;    16'd49589: out <= 16'h037B;    16'd49590: out <= 16'h0AF3;    16'd49591: out <= 16'h05EB;
    16'd49592: out <= 16'h08B8;    16'd49593: out <= 16'h06B4;    16'd49594: out <= 16'h08A6;    16'd49595: out <= 16'hFC80;
    16'd49596: out <= 16'hFFCB;    16'd49597: out <= 16'h089D;    16'd49598: out <= 16'h05A8;    16'd49599: out <= 16'h09F8;
    16'd49600: out <= 16'h09B6;    16'd49601: out <= 16'hFF31;    16'd49602: out <= 16'h0515;    16'd49603: out <= 16'h0069;
    16'd49604: out <= 16'h0393;    16'd49605: out <= 16'h0268;    16'd49606: out <= 16'hFF11;    16'd49607: out <= 16'h023B;
    16'd49608: out <= 16'hFE8E;    16'd49609: out <= 16'hFEEA;    16'd49610: out <= 16'h027E;    16'd49611: out <= 16'hFF0C;
    16'd49612: out <= 16'hFD78;    16'd49613: out <= 16'hFF11;    16'd49614: out <= 16'hFC88;    16'd49615: out <= 16'h0541;
    16'd49616: out <= 16'h06BB;    16'd49617: out <= 16'hFEA6;    16'd49618: out <= 16'hFC49;    16'd49619: out <= 16'h0134;
    16'd49620: out <= 16'hFA33;    16'd49621: out <= 16'hFE5C;    16'd49622: out <= 16'h02E1;    16'd49623: out <= 16'hFA15;
    16'd49624: out <= 16'hFCBA;    16'd49625: out <= 16'h00DA;    16'd49626: out <= 16'hFF52;    16'd49627: out <= 16'h0353;
    16'd49628: out <= 16'hFEF1;    16'd49629: out <= 16'h046C;    16'd49630: out <= 16'h0B4F;    16'd49631: out <= 16'h04CF;
    16'd49632: out <= 16'hFDA4;    16'd49633: out <= 16'h0205;    16'd49634: out <= 16'h022A;    16'd49635: out <= 16'h00F7;
    16'd49636: out <= 16'hFCCB;    16'd49637: out <= 16'hFF05;    16'd49638: out <= 16'h06CB;    16'd49639: out <= 16'h08ED;
    16'd49640: out <= 16'h01FE;    16'd49641: out <= 16'h08A9;    16'd49642: out <= 16'h007C;    16'd49643: out <= 16'hFA97;
    16'd49644: out <= 16'h01A7;    16'd49645: out <= 16'h05E3;    16'd49646: out <= 16'h0160;    16'd49647: out <= 16'h0521;
    16'd49648: out <= 16'hFE33;    16'd49649: out <= 16'hF915;    16'd49650: out <= 16'hFD4C;    16'd49651: out <= 16'hF9DA;
    16'd49652: out <= 16'hF7B9;    16'd49653: out <= 16'hFEB9;    16'd49654: out <= 16'hFA78;    16'd49655: out <= 16'h03CF;
    16'd49656: out <= 16'hFEA7;    16'd49657: out <= 16'h00DC;    16'd49658: out <= 16'h01AB;    16'd49659: out <= 16'h02D7;
    16'd49660: out <= 16'hFC39;    16'd49661: out <= 16'hFEA0;    16'd49662: out <= 16'hFF6E;    16'd49663: out <= 16'hFF2D;
    16'd49664: out <= 16'h0402;    16'd49665: out <= 16'h0102;    16'd49666: out <= 16'hFC36;    16'd49667: out <= 16'hF7C2;
    16'd49668: out <= 16'h0064;    16'd49669: out <= 16'h060C;    16'd49670: out <= 16'hF8DD;    16'd49671: out <= 16'h0352;
    16'd49672: out <= 16'h009D;    16'd49673: out <= 16'hFF94;    16'd49674: out <= 16'h00E3;    16'd49675: out <= 16'hFCF4;
    16'd49676: out <= 16'hFB42;    16'd49677: out <= 16'h056E;    16'd49678: out <= 16'hFCB3;    16'd49679: out <= 16'h0053;
    16'd49680: out <= 16'h00BD;    16'd49681: out <= 16'h0363;    16'd49682: out <= 16'h0885;    16'd49683: out <= 16'h0301;
    16'd49684: out <= 16'hFF51;    16'd49685: out <= 16'h02EB;    16'd49686: out <= 16'hFD50;    16'd49687: out <= 16'h0026;
    16'd49688: out <= 16'hFD9A;    16'd49689: out <= 16'hFC1D;    16'd49690: out <= 16'hFDF4;    16'd49691: out <= 16'hFDB0;
    16'd49692: out <= 16'hF6DD;    16'd49693: out <= 16'h0365;    16'd49694: out <= 16'hF657;    16'd49695: out <= 16'hFECF;
    16'd49696: out <= 16'hFF72;    16'd49697: out <= 16'hFE9A;    16'd49698: out <= 16'hFF08;    16'd49699: out <= 16'h03A8;
    16'd49700: out <= 16'h03D1;    16'd49701: out <= 16'h0496;    16'd49702: out <= 16'h0007;    16'd49703: out <= 16'hFEC8;
    16'd49704: out <= 16'hFF40;    16'd49705: out <= 16'h02DC;    16'd49706: out <= 16'hFAF3;    16'd49707: out <= 16'h0381;
    16'd49708: out <= 16'h08BE;    16'd49709: out <= 16'h0155;    16'd49710: out <= 16'h0800;    16'd49711: out <= 16'h0737;
    16'd49712: out <= 16'hFE2D;    16'd49713: out <= 16'h0F58;    16'd49714: out <= 16'hFB4C;    16'd49715: out <= 16'hFEA8;
    16'd49716: out <= 16'h057B;    16'd49717: out <= 16'h06D7;    16'd49718: out <= 16'h05C4;    16'd49719: out <= 16'h04F4;
    16'd49720: out <= 16'h0987;    16'd49721: out <= 16'h00D3;    16'd49722: out <= 16'h036D;    16'd49723: out <= 16'h0691;
    16'd49724: out <= 16'h0A1B;    16'd49725: out <= 16'h0310;    16'd49726: out <= 16'hFF8D;    16'd49727: out <= 16'h0308;
    16'd49728: out <= 16'h0228;    16'd49729: out <= 16'h053A;    16'd49730: out <= 16'h02DB;    16'd49731: out <= 16'hFF3D;
    16'd49732: out <= 16'h0204;    16'd49733: out <= 16'h08A9;    16'd49734: out <= 16'h02DB;    16'd49735: out <= 16'h06AE;
    16'd49736: out <= 16'h0194;    16'd49737: out <= 16'h04ED;    16'd49738: out <= 16'h0386;    16'd49739: out <= 16'h054F;
    16'd49740: out <= 16'h0181;    16'd49741: out <= 16'h045B;    16'd49742: out <= 16'h0BC3;    16'd49743: out <= 16'hFBC7;
    16'd49744: out <= 16'hFF78;    16'd49745: out <= 16'h083A;    16'd49746: out <= 16'hFE1B;    16'd49747: out <= 16'hFF45;
    16'd49748: out <= 16'h03BE;    16'd49749: out <= 16'h03F5;    16'd49750: out <= 16'hFCDC;    16'd49751: out <= 16'h080A;
    16'd49752: out <= 16'h03FA;    16'd49753: out <= 16'h02D7;    16'd49754: out <= 16'hFC24;    16'd49755: out <= 16'h0568;
    16'd49756: out <= 16'hFACE;    16'd49757: out <= 16'h0268;    16'd49758: out <= 16'h0168;    16'd49759: out <= 16'h0615;
    16'd49760: out <= 16'h055B;    16'd49761: out <= 16'h011F;    16'd49762: out <= 16'h067B;    16'd49763: out <= 16'hFFD9;
    16'd49764: out <= 16'h051E;    16'd49765: out <= 16'h015F;    16'd49766: out <= 16'h00C1;    16'd49767: out <= 16'h062C;
    16'd49768: out <= 16'h03F7;    16'd49769: out <= 16'hFFE7;    16'd49770: out <= 16'h0BD7;    16'd49771: out <= 16'h02CB;
    16'd49772: out <= 16'hFDA0;    16'd49773: out <= 16'h0CD6;    16'd49774: out <= 16'h05A3;    16'd49775: out <= 16'h0912;
    16'd49776: out <= 16'h036A;    16'd49777: out <= 16'h0B7D;    16'd49778: out <= 16'h0534;    16'd49779: out <= 16'hFCFD;
    16'd49780: out <= 16'h05C7;    16'd49781: out <= 16'h052E;    16'd49782: out <= 16'h0777;    16'd49783: out <= 16'h0751;
    16'd49784: out <= 16'h020F;    16'd49785: out <= 16'h069B;    16'd49786: out <= 16'h01F9;    16'd49787: out <= 16'h010B;
    16'd49788: out <= 16'h05F2;    16'd49789: out <= 16'h0398;    16'd49790: out <= 16'h022F;    16'd49791: out <= 16'h00BD;
    16'd49792: out <= 16'h061F;    16'd49793: out <= 16'h0709;    16'd49794: out <= 16'h075B;    16'd49795: out <= 16'h08AA;
    16'd49796: out <= 16'h03FB;    16'd49797: out <= 16'h06FA;    16'd49798: out <= 16'h0105;    16'd49799: out <= 16'h03F8;
    16'd49800: out <= 16'h040F;    16'd49801: out <= 16'hFF47;    16'd49802: out <= 16'h01A5;    16'd49803: out <= 16'h01B5;
    16'd49804: out <= 16'h0046;    16'd49805: out <= 16'h013A;    16'd49806: out <= 16'hFFBD;    16'd49807: out <= 16'h0510;
    16'd49808: out <= 16'h0C66;    16'd49809: out <= 16'h02F6;    16'd49810: out <= 16'hFFF5;    16'd49811: out <= 16'hFCEB;
    16'd49812: out <= 16'h013A;    16'd49813: out <= 16'h02BA;    16'd49814: out <= 16'h059E;    16'd49815: out <= 16'h096C;
    16'd49816: out <= 16'h015B;    16'd49817: out <= 16'h0227;    16'd49818: out <= 16'h0082;    16'd49819: out <= 16'h0311;
    16'd49820: out <= 16'h059E;    16'd49821: out <= 16'h0778;    16'd49822: out <= 16'h08FE;    16'd49823: out <= 16'h0643;
    16'd49824: out <= 16'h091F;    16'd49825: out <= 16'h0290;    16'd49826: out <= 16'h0319;    16'd49827: out <= 16'h0516;
    16'd49828: out <= 16'h033D;    16'd49829: out <= 16'h0434;    16'd49830: out <= 16'h035C;    16'd49831: out <= 16'h0477;
    16'd49832: out <= 16'hF9A5;    16'd49833: out <= 16'h083B;    16'd49834: out <= 16'h046B;    16'd49835: out <= 16'h0A9F;
    16'd49836: out <= 16'h062B;    16'd49837: out <= 16'h02F2;    16'd49838: out <= 16'h0202;    16'd49839: out <= 16'h0395;
    16'd49840: out <= 16'h0623;    16'd49841: out <= 16'h069F;    16'd49842: out <= 16'h09FC;    16'd49843: out <= 16'h02E8;
    16'd49844: out <= 16'h00CE;    16'd49845: out <= 16'hF9AE;    16'd49846: out <= 16'h045D;    16'd49847: out <= 16'h005B;
    16'd49848: out <= 16'h03E0;    16'd49849: out <= 16'h080F;    16'd49850: out <= 16'h0269;    16'd49851: out <= 16'h058D;
    16'd49852: out <= 16'h05BB;    16'd49853: out <= 16'h043A;    16'd49854: out <= 16'h0865;    16'd49855: out <= 16'h0432;
    16'd49856: out <= 16'hFD83;    16'd49857: out <= 16'h04E7;    16'd49858: out <= 16'h05E2;    16'd49859: out <= 16'h0583;
    16'd49860: out <= 16'h00B2;    16'd49861: out <= 16'h03E2;    16'd49862: out <= 16'hFC2F;    16'd49863: out <= 16'hFF65;
    16'd49864: out <= 16'h021B;    16'd49865: out <= 16'h00C7;    16'd49866: out <= 16'h0A78;    16'd49867: out <= 16'hFFC9;
    16'd49868: out <= 16'h03C6;    16'd49869: out <= 16'h06E3;    16'd49870: out <= 16'h00BA;    16'd49871: out <= 16'h01BE;
    16'd49872: out <= 16'hF819;    16'd49873: out <= 16'h0142;    16'd49874: out <= 16'hFF3B;    16'd49875: out <= 16'h006E;
    16'd49876: out <= 16'h03C1;    16'd49877: out <= 16'h018B;    16'd49878: out <= 16'hFFC5;    16'd49879: out <= 16'hFC86;
    16'd49880: out <= 16'h038D;    16'd49881: out <= 16'h02E7;    16'd49882: out <= 16'hFF0B;    16'd49883: out <= 16'h0417;
    16'd49884: out <= 16'h035E;    16'd49885: out <= 16'hFF60;    16'd49886: out <= 16'hFEC4;    16'd49887: out <= 16'hFE88;
    16'd49888: out <= 16'hFAB8;    16'd49889: out <= 16'hFC73;    16'd49890: out <= 16'h02DF;    16'd49891: out <= 16'h0932;
    16'd49892: out <= 16'hF61E;    16'd49893: out <= 16'h0020;    16'd49894: out <= 16'hFBC0;    16'd49895: out <= 16'hFABB;
    16'd49896: out <= 16'hFAEA;    16'd49897: out <= 16'hFFC3;    16'd49898: out <= 16'hFBBF;    16'd49899: out <= 16'hFD4F;
    16'd49900: out <= 16'h0083;    16'd49901: out <= 16'hFA78;    16'd49902: out <= 16'hFF98;    16'd49903: out <= 16'hFF2A;
    16'd49904: out <= 16'hFD4D;    16'd49905: out <= 16'h0768;    16'd49906: out <= 16'hFF50;    16'd49907: out <= 16'hFEA9;
    16'd49908: out <= 16'h0165;    16'd49909: out <= 16'hFAC0;    16'd49910: out <= 16'h026B;    16'd49911: out <= 16'hFB51;
    16'd49912: out <= 16'h07E4;    16'd49913: out <= 16'h022A;    16'd49914: out <= 16'hFAA3;    16'd49915: out <= 16'hFED9;
    16'd49916: out <= 16'h0335;    16'd49917: out <= 16'hFE87;    16'd49918: out <= 16'hFBF6;    16'd49919: out <= 16'h013C;
    16'd49920: out <= 16'h02FA;    16'd49921: out <= 16'h0581;    16'd49922: out <= 16'hF7EB;    16'd49923: out <= 16'h03CC;
    16'd49924: out <= 16'h0772;    16'd49925: out <= 16'h049D;    16'd49926: out <= 16'h0332;    16'd49927: out <= 16'hFDA5;
    16'd49928: out <= 16'h019F;    16'd49929: out <= 16'hFEE4;    16'd49930: out <= 16'h024D;    16'd49931: out <= 16'h04AE;
    16'd49932: out <= 16'h0019;    16'd49933: out <= 16'h0332;    16'd49934: out <= 16'hFF4D;    16'd49935: out <= 16'hFC03;
    16'd49936: out <= 16'h03F2;    16'd49937: out <= 16'h0040;    16'd49938: out <= 16'hFD7A;    16'd49939: out <= 16'h0169;
    16'd49940: out <= 16'hFD1F;    16'd49941: out <= 16'h0476;    16'd49942: out <= 16'h03EE;    16'd49943: out <= 16'hFA6A;
    16'd49944: out <= 16'h002E;    16'd49945: out <= 16'h03E1;    16'd49946: out <= 16'hFA47;    16'd49947: out <= 16'h03FE;
    16'd49948: out <= 16'hFA91;    16'd49949: out <= 16'h0625;    16'd49950: out <= 16'h05E5;    16'd49951: out <= 16'hFAFC;
    16'd49952: out <= 16'hFC9F;    16'd49953: out <= 16'h03BF;    16'd49954: out <= 16'hFC6C;    16'd49955: out <= 16'h0742;
    16'd49956: out <= 16'hFE17;    16'd49957: out <= 16'hFF53;    16'd49958: out <= 16'hFFF1;    16'd49959: out <= 16'hFF9B;
    16'd49960: out <= 16'hFF6D;    16'd49961: out <= 16'h02D7;    16'd49962: out <= 16'h0374;    16'd49963: out <= 16'h03EB;
    16'd49964: out <= 16'h03B5;    16'd49965: out <= 16'h06B9;    16'd49966: out <= 16'h0BAB;    16'd49967: out <= 16'hFE26;
    16'd49968: out <= 16'h0CDF;    16'd49969: out <= 16'h0618;    16'd49970: out <= 16'hFC7E;    16'd49971: out <= 16'h0357;
    16'd49972: out <= 16'h0130;    16'd49973: out <= 16'h036E;    16'd49974: out <= 16'h0421;    16'd49975: out <= 16'h007F;
    16'd49976: out <= 16'h01C1;    16'd49977: out <= 16'h0983;    16'd49978: out <= 16'h0487;    16'd49979: out <= 16'h05FC;
    16'd49980: out <= 16'h03B3;    16'd49981: out <= 16'h0573;    16'd49982: out <= 16'h06A0;    16'd49983: out <= 16'hFF1A;
    16'd49984: out <= 16'h00DD;    16'd49985: out <= 16'h0628;    16'd49986: out <= 16'h01B4;    16'd49987: out <= 16'hFB1A;
    16'd49988: out <= 16'h0640;    16'd49989: out <= 16'h0874;    16'd49990: out <= 16'h0406;    16'd49991: out <= 16'h0886;
    16'd49992: out <= 16'h0452;    16'd49993: out <= 16'h0979;    16'd49994: out <= 16'h0366;    16'd49995: out <= 16'h0440;
    16'd49996: out <= 16'h063E;    16'd49997: out <= 16'h01DE;    16'd49998: out <= 16'h00CF;    16'd49999: out <= 16'h00E0;
    16'd50000: out <= 16'hFF6B;    16'd50001: out <= 16'h06A6;    16'd50002: out <= 16'h0BFC;    16'd50003: out <= 16'h0368;
    16'd50004: out <= 16'h027B;    16'd50005: out <= 16'hFE56;    16'd50006: out <= 16'h0730;    16'd50007: out <= 16'hFF40;
    16'd50008: out <= 16'h01F7;    16'd50009: out <= 16'h019C;    16'd50010: out <= 16'h08D0;    16'd50011: out <= 16'h096A;
    16'd50012: out <= 16'h06ED;    16'd50013: out <= 16'hFD7E;    16'd50014: out <= 16'h0605;    16'd50015: out <= 16'h0A2F;
    16'd50016: out <= 16'h0516;    16'd50017: out <= 16'h063E;    16'd50018: out <= 16'hFD6A;    16'd50019: out <= 16'h0038;
    16'd50020: out <= 16'h006F;    16'd50021: out <= 16'h03D0;    16'd50022: out <= 16'hFFDF;    16'd50023: out <= 16'h006A;
    16'd50024: out <= 16'h040C;    16'd50025: out <= 16'h07AF;    16'd50026: out <= 16'h03DE;    16'd50027: out <= 16'hFE29;
    16'd50028: out <= 16'h0A1E;    16'd50029: out <= 16'h04A0;    16'd50030: out <= 16'h06B9;    16'd50031: out <= 16'h08E6;
    16'd50032: out <= 16'h02EF;    16'd50033: out <= 16'h022C;    16'd50034: out <= 16'h0715;    16'd50035: out <= 16'hFED2;
    16'd50036: out <= 16'h0765;    16'd50037: out <= 16'h093C;    16'd50038: out <= 16'h057E;    16'd50039: out <= 16'h0733;
    16'd50040: out <= 16'h067E;    16'd50041: out <= 16'hFF33;    16'd50042: out <= 16'h0828;    16'd50043: out <= 16'h035F;
    16'd50044: out <= 16'h032E;    16'd50045: out <= 16'h04F3;    16'd50046: out <= 16'h012D;    16'd50047: out <= 16'h0411;
    16'd50048: out <= 16'h0717;    16'd50049: out <= 16'h02C7;    16'd50050: out <= 16'h0593;    16'd50051: out <= 16'h0687;
    16'd50052: out <= 16'hFFE4;    16'd50053: out <= 16'h0973;    16'd50054: out <= 16'h05F3;    16'd50055: out <= 16'h039F;
    16'd50056: out <= 16'h074C;    16'd50057: out <= 16'h0504;    16'd50058: out <= 16'h03C4;    16'd50059: out <= 16'h07F3;
    16'd50060: out <= 16'h0241;    16'd50061: out <= 16'h04D6;    16'd50062: out <= 16'h0648;    16'd50063: out <= 16'h04E2;
    16'd50064: out <= 16'h050D;    16'd50065: out <= 16'h0315;    16'd50066: out <= 16'h050D;    16'd50067: out <= 16'h08FE;
    16'd50068: out <= 16'h01F1;    16'd50069: out <= 16'hFB27;    16'd50070: out <= 16'h0745;    16'd50071: out <= 16'h0AB9;
    16'd50072: out <= 16'h08F1;    16'd50073: out <= 16'h0CE3;    16'd50074: out <= 16'h01A0;    16'd50075: out <= 16'h089B;
    16'd50076: out <= 16'hFC18;    16'd50077: out <= 16'h0402;    16'd50078: out <= 16'h0182;    16'd50079: out <= 16'h0350;
    16'd50080: out <= 16'h07C7;    16'd50081: out <= 16'h0734;    16'd50082: out <= 16'h08E6;    16'd50083: out <= 16'hFE4D;
    16'd50084: out <= 16'h04D3;    16'd50085: out <= 16'h0109;    16'd50086: out <= 16'h00E5;    16'd50087: out <= 16'h0243;
    16'd50088: out <= 16'h021D;    16'd50089: out <= 16'hFFC0;    16'd50090: out <= 16'h0A21;    16'd50091: out <= 16'h0800;
    16'd50092: out <= 16'h055E;    16'd50093: out <= 16'h05A4;    16'd50094: out <= 16'h07C2;    16'd50095: out <= 16'h0150;
    16'd50096: out <= 16'h000E;    16'd50097: out <= 16'h04A3;    16'd50098: out <= 16'h08D0;    16'd50099: out <= 16'h0619;
    16'd50100: out <= 16'h06D2;    16'd50101: out <= 16'h038D;    16'd50102: out <= 16'h0859;    16'd50103: out <= 16'h092F;
    16'd50104: out <= 16'h05B0;    16'd50105: out <= 16'h05E7;    16'd50106: out <= 16'h09E2;    16'd50107: out <= 16'h0586;
    16'd50108: out <= 16'h01E1;    16'd50109: out <= 16'h060F;    16'd50110: out <= 16'hFFE5;    16'd50111: out <= 16'h08F8;
    16'd50112: out <= 16'hFCA6;    16'd50113: out <= 16'h083D;    16'd50114: out <= 16'hFF4E;    16'd50115: out <= 16'h0287;
    16'd50116: out <= 16'h0369;    16'd50117: out <= 16'hFB24;    16'd50118: out <= 16'h01C4;    16'd50119: out <= 16'hFEA4;
    16'd50120: out <= 16'h0398;    16'd50121: out <= 16'hF95F;    16'd50122: out <= 16'hF67A;    16'd50123: out <= 16'hFE01;
    16'd50124: out <= 16'h011F;    16'd50125: out <= 16'hFCF1;    16'd50126: out <= 16'hF9B6;    16'd50127: out <= 16'hFE10;
    16'd50128: out <= 16'hFFDA;    16'd50129: out <= 16'hFAB7;    16'd50130: out <= 16'hFEF5;    16'd50131: out <= 16'h066B;
    16'd50132: out <= 16'hFE2D;    16'd50133: out <= 16'h0118;    16'd50134: out <= 16'h09A6;    16'd50135: out <= 16'hFF5D;
    16'd50136: out <= 16'hFA8D;    16'd50137: out <= 16'hFD55;    16'd50138: out <= 16'hFDC3;    16'd50139: out <= 16'hF939;
    16'd50140: out <= 16'hFD04;    16'd50141: out <= 16'h02AB;    16'd50142: out <= 16'hFECE;    16'd50143: out <= 16'hFE2D;
    16'd50144: out <= 16'hFDDD;    16'd50145: out <= 16'hFCCF;    16'd50146: out <= 16'hFB7B;    16'd50147: out <= 16'hFD04;
    16'd50148: out <= 16'hFDC8;    16'd50149: out <= 16'h03E1;    16'd50150: out <= 16'h0102;    16'd50151: out <= 16'hF5AF;
    16'd50152: out <= 16'h04A0;    16'd50153: out <= 16'h0504;    16'd50154: out <= 16'h00C9;    16'd50155: out <= 16'hF2BD;
    16'd50156: out <= 16'h02AC;    16'd50157: out <= 16'hFC81;    16'd50158: out <= 16'hFD7A;    16'd50159: out <= 16'hFB7C;
    16'd50160: out <= 16'hFF0B;    16'd50161: out <= 16'hFE0E;    16'd50162: out <= 16'h01DF;    16'd50163: out <= 16'hFF4A;
    16'd50164: out <= 16'hFF41;    16'd50165: out <= 16'h023B;    16'd50166: out <= 16'h06C8;    16'd50167: out <= 16'h04E6;
    16'd50168: out <= 16'h0510;    16'd50169: out <= 16'h04C3;    16'd50170: out <= 16'hFD2A;    16'd50171: out <= 16'h0024;
    16'd50172: out <= 16'h0007;    16'd50173: out <= 16'hFF8A;    16'd50174: out <= 16'hFE06;    16'd50175: out <= 16'hFFD4;
    16'd50176: out <= 16'h006C;    16'd50177: out <= 16'hFF6F;    16'd50178: out <= 16'h05E4;    16'd50179: out <= 16'hFCA9;
    16'd50180: out <= 16'h01F9;    16'd50181: out <= 16'hFE00;    16'd50182: out <= 16'hFDD9;    16'd50183: out <= 16'h014D;
    16'd50184: out <= 16'h021A;    16'd50185: out <= 16'h030B;    16'd50186: out <= 16'hFBE3;    16'd50187: out <= 16'h0051;
    16'd50188: out <= 16'hFF86;    16'd50189: out <= 16'hFF40;    16'd50190: out <= 16'hFCD2;    16'd50191: out <= 16'h0555;
    16'd50192: out <= 16'hFF18;    16'd50193: out <= 16'h00A9;    16'd50194: out <= 16'hFF6F;    16'd50195: out <= 16'hFE01;
    16'd50196: out <= 16'h01A3;    16'd50197: out <= 16'h06D3;    16'd50198: out <= 16'h050B;    16'd50199: out <= 16'hFBC6;
    16'd50200: out <= 16'h01CF;    16'd50201: out <= 16'h025A;    16'd50202: out <= 16'hFE57;    16'd50203: out <= 16'h0266;
    16'd50204: out <= 16'h06A4;    16'd50205: out <= 16'h0154;    16'd50206: out <= 16'hFC16;    16'd50207: out <= 16'h0559;
    16'd50208: out <= 16'h04C7;    16'd50209: out <= 16'hFF38;    16'd50210: out <= 16'hFF19;    16'd50211: out <= 16'h040B;
    16'd50212: out <= 16'hFED4;    16'd50213: out <= 16'h0546;    16'd50214: out <= 16'h008E;    16'd50215: out <= 16'h0050;
    16'd50216: out <= 16'h0642;    16'd50217: out <= 16'h0115;    16'd50218: out <= 16'h045D;    16'd50219: out <= 16'h046E;
    16'd50220: out <= 16'h016D;    16'd50221: out <= 16'h01D4;    16'd50222: out <= 16'h0298;    16'd50223: out <= 16'hFFBA;
    16'd50224: out <= 16'hFB2C;    16'd50225: out <= 16'h0604;    16'd50226: out <= 16'hFF15;    16'd50227: out <= 16'h04C4;
    16'd50228: out <= 16'h055F;    16'd50229: out <= 16'h0448;    16'd50230: out <= 16'h0404;    16'd50231: out <= 16'hFE1F;
    16'd50232: out <= 16'h0212;    16'd50233: out <= 16'h03B8;    16'd50234: out <= 16'hFBD7;    16'd50235: out <= 16'h057D;
    16'd50236: out <= 16'h02F1;    16'd50237: out <= 16'hFF5B;    16'd50238: out <= 16'h080A;    16'd50239: out <= 16'h008F;
    16'd50240: out <= 16'h05B4;    16'd50241: out <= 16'h030C;    16'd50242: out <= 16'hFDAC;    16'd50243: out <= 16'h06E2;
    16'd50244: out <= 16'h055B;    16'd50245: out <= 16'hFD74;    16'd50246: out <= 16'h0572;    16'd50247: out <= 16'h0052;
    16'd50248: out <= 16'h08C9;    16'd50249: out <= 16'h091E;    16'd50250: out <= 16'h07C0;    16'd50251: out <= 16'h038E;
    16'd50252: out <= 16'h009F;    16'd50253: out <= 16'hFDA2;    16'd50254: out <= 16'h089F;    16'd50255: out <= 16'h07BA;
    16'd50256: out <= 16'h08C9;    16'd50257: out <= 16'h0AC4;    16'd50258: out <= 16'h05F5;    16'd50259: out <= 16'h05D3;
    16'd50260: out <= 16'h086E;    16'd50261: out <= 16'h085B;    16'd50262: out <= 16'h0609;    16'd50263: out <= 16'hFFA8;
    16'd50264: out <= 16'h0700;    16'd50265: out <= 16'h0580;    16'd50266: out <= 16'h009B;    16'd50267: out <= 16'h0266;
    16'd50268: out <= 16'h0384;    16'd50269: out <= 16'hFE9D;    16'd50270: out <= 16'h0522;    16'd50271: out <= 16'h0711;
    16'd50272: out <= 16'h0684;    16'd50273: out <= 16'hFF3C;    16'd50274: out <= 16'h09D5;    16'd50275: out <= 16'h0383;
    16'd50276: out <= 16'h052E;    16'd50277: out <= 16'h0497;    16'd50278: out <= 16'hFD30;    16'd50279: out <= 16'h0566;
    16'd50280: out <= 16'h004D;    16'd50281: out <= 16'h0882;    16'd50282: out <= 16'h04A1;    16'd50283: out <= 16'hFC6F;
    16'd50284: out <= 16'h054B;    16'd50285: out <= 16'hFE68;    16'd50286: out <= 16'hFD0A;    16'd50287: out <= 16'h01E5;
    16'd50288: out <= 16'h0012;    16'd50289: out <= 16'h0347;    16'd50290: out <= 16'h02C2;    16'd50291: out <= 16'h03E4;
    16'd50292: out <= 16'hFCAE;    16'd50293: out <= 16'h07AE;    16'd50294: out <= 16'hFD40;    16'd50295: out <= 16'hFC03;
    16'd50296: out <= 16'hFF70;    16'd50297: out <= 16'h0413;    16'd50298: out <= 16'h05BD;    16'd50299: out <= 16'h062F;
    16'd50300: out <= 16'h0763;    16'd50301: out <= 16'h01AF;    16'd50302: out <= 16'h002A;    16'd50303: out <= 16'h09EB;
    16'd50304: out <= 16'h007E;    16'd50305: out <= 16'h0229;    16'd50306: out <= 16'h03CD;    16'd50307: out <= 16'h07F7;
    16'd50308: out <= 16'h02BD;    16'd50309: out <= 16'h0700;    16'd50310: out <= 16'h032C;    16'd50311: out <= 16'hFF5B;
    16'd50312: out <= 16'h037B;    16'd50313: out <= 16'h080D;    16'd50314: out <= 16'h0408;    16'd50315: out <= 16'h02DE;
    16'd50316: out <= 16'h04FB;    16'd50317: out <= 16'h05D5;    16'd50318: out <= 16'h006B;    16'd50319: out <= 16'h02B3;
    16'd50320: out <= 16'h09BC;    16'd50321: out <= 16'h03EA;    16'd50322: out <= 16'h0509;    16'd50323: out <= 16'h0366;
    16'd50324: out <= 16'hFE1E;    16'd50325: out <= 16'h01BD;    16'd50326: out <= 16'h00ED;    16'd50327: out <= 16'h061B;
    16'd50328: out <= 16'h038A;    16'd50329: out <= 16'hF929;    16'd50330: out <= 16'h0201;    16'd50331: out <= 16'h0396;
    16'd50332: out <= 16'h01BB;    16'd50333: out <= 16'h05C4;    16'd50334: out <= 16'hFED9;    16'd50335: out <= 16'h0539;
    16'd50336: out <= 16'h0621;    16'd50337: out <= 16'h0881;    16'd50338: out <= 16'h059F;    16'd50339: out <= 16'h00CD;
    16'd50340: out <= 16'h04A7;    16'd50341: out <= 16'h0122;    16'd50342: out <= 16'h015D;    16'd50343: out <= 16'h05BA;
    16'd50344: out <= 16'h03E0;    16'd50345: out <= 16'h0325;    16'd50346: out <= 16'h0774;    16'd50347: out <= 16'h0972;
    16'd50348: out <= 16'h04B0;    16'd50349: out <= 16'hFC76;    16'd50350: out <= 16'h0552;    16'd50351: out <= 16'h097E;
    16'd50352: out <= 16'h03CE;    16'd50353: out <= 16'h0449;    16'd50354: out <= 16'h0866;    16'd50355: out <= 16'h02CE;
    16'd50356: out <= 16'h0813;    16'd50357: out <= 16'hFFEC;    16'd50358: out <= 16'h00E8;    16'd50359: out <= 16'h07C8;
    16'd50360: out <= 16'h0A18;    16'd50361: out <= 16'hFEAA;    16'd50362: out <= 16'h0468;    16'd50363: out <= 16'h03B2;
    16'd50364: out <= 16'h0A07;    16'd50365: out <= 16'h01DA;    16'd50366: out <= 16'h07A5;    16'd50367: out <= 16'h0399;
    16'd50368: out <= 16'h0938;    16'd50369: out <= 16'h0774;    16'd50370: out <= 16'h0876;    16'd50371: out <= 16'h0056;
    16'd50372: out <= 16'hF7C9;    16'd50373: out <= 16'hFE91;    16'd50374: out <= 16'hFE83;    16'd50375: out <= 16'h0396;
    16'd50376: out <= 16'h01C3;    16'd50377: out <= 16'h0A44;    16'd50378: out <= 16'hFD24;    16'd50379: out <= 16'h010A;
    16'd50380: out <= 16'h0472;    16'd50381: out <= 16'h00A0;    16'd50382: out <= 16'h00EA;    16'd50383: out <= 16'h0046;
    16'd50384: out <= 16'h041A;    16'd50385: out <= 16'h01D2;    16'd50386: out <= 16'h0268;    16'd50387: out <= 16'hFEBB;
    16'd50388: out <= 16'h008F;    16'd50389: out <= 16'hFC22;    16'd50390: out <= 16'h0246;    16'd50391: out <= 16'hF8A3;
    16'd50392: out <= 16'h01D2;    16'd50393: out <= 16'hFF0C;    16'd50394: out <= 16'hFC44;    16'd50395: out <= 16'hFD4C;
    16'd50396: out <= 16'hFF2F;    16'd50397: out <= 16'hFC29;    16'd50398: out <= 16'hFE47;    16'd50399: out <= 16'hFD91;
    16'd50400: out <= 16'hF9FE;    16'd50401: out <= 16'h02FD;    16'd50402: out <= 16'h037C;    16'd50403: out <= 16'hFAA8;
    16'd50404: out <= 16'hFE4E;    16'd50405: out <= 16'h00F5;    16'd50406: out <= 16'hFE54;    16'd50407: out <= 16'h03DF;
    16'd50408: out <= 16'h070C;    16'd50409: out <= 16'h016A;    16'd50410: out <= 16'hFBCD;    16'd50411: out <= 16'hFF61;
    16'd50412: out <= 16'h01DC;    16'd50413: out <= 16'hFF71;    16'd50414: out <= 16'hFADF;    16'd50415: out <= 16'h0480;
    16'd50416: out <= 16'hFA85;    16'd50417: out <= 16'hFA89;    16'd50418: out <= 16'h00E7;    16'd50419: out <= 16'hFBDC;
    16'd50420: out <= 16'h0338;    16'd50421: out <= 16'h0192;    16'd50422: out <= 16'h039A;    16'd50423: out <= 16'hFDF0;
    16'd50424: out <= 16'h025E;    16'd50425: out <= 16'h03BA;    16'd50426: out <= 16'hF80C;    16'd50427: out <= 16'h0190;
    16'd50428: out <= 16'h002A;    16'd50429: out <= 16'h020A;    16'd50430: out <= 16'h0285;    16'd50431: out <= 16'hFBB3;
    16'd50432: out <= 16'h01E9;    16'd50433: out <= 16'h0463;    16'd50434: out <= 16'h023F;    16'd50435: out <= 16'hFC45;
    16'd50436: out <= 16'h020E;    16'd50437: out <= 16'h07E6;    16'd50438: out <= 16'h015A;    16'd50439: out <= 16'h05B3;
    16'd50440: out <= 16'hFA3A;    16'd50441: out <= 16'h01A9;    16'd50442: out <= 16'h0326;    16'd50443: out <= 16'h029D;
    16'd50444: out <= 16'h02A6;    16'd50445: out <= 16'h034D;    16'd50446: out <= 16'hFC4C;    16'd50447: out <= 16'hFC9E;
    16'd50448: out <= 16'hFFC3;    16'd50449: out <= 16'h01AA;    16'd50450: out <= 16'h01A5;    16'd50451: out <= 16'hFF47;
    16'd50452: out <= 16'hFE67;    16'd50453: out <= 16'hFDCE;    16'd50454: out <= 16'h01AC;    16'd50455: out <= 16'h05CE;
    16'd50456: out <= 16'h0610;    16'd50457: out <= 16'h0673;    16'd50458: out <= 16'hFE85;    16'd50459: out <= 16'h026E;
    16'd50460: out <= 16'h0275;    16'd50461: out <= 16'hFF35;    16'd50462: out <= 16'h011D;    16'd50463: out <= 16'hFC05;
    16'd50464: out <= 16'hFA8B;    16'd50465: out <= 16'hFBA7;    16'd50466: out <= 16'h03FD;    16'd50467: out <= 16'hFD07;
    16'd50468: out <= 16'h006A;    16'd50469: out <= 16'hFDA2;    16'd50470: out <= 16'h03EE;    16'd50471: out <= 16'h0240;
    16'd50472: out <= 16'h03C6;    16'd50473: out <= 16'h05E0;    16'd50474: out <= 16'h01A5;    16'd50475: out <= 16'h02D9;
    16'd50476: out <= 16'h041B;    16'd50477: out <= 16'h0222;    16'd50478: out <= 16'h0D27;    16'd50479: out <= 16'h0B1F;
    16'd50480: out <= 16'hFCA3;    16'd50481: out <= 16'h0593;    16'd50482: out <= 16'hFDD1;    16'd50483: out <= 16'h05D5;
    16'd50484: out <= 16'h0526;    16'd50485: out <= 16'h001F;    16'd50486: out <= 16'h0B1A;    16'd50487: out <= 16'h0231;
    16'd50488: out <= 16'h05CA;    16'd50489: out <= 16'h03ED;    16'd50490: out <= 16'h04FB;    16'd50491: out <= 16'h0739;
    16'd50492: out <= 16'h02F5;    16'd50493: out <= 16'h0213;    16'd50494: out <= 16'h02C9;    16'd50495: out <= 16'h0474;
    16'd50496: out <= 16'h065A;    16'd50497: out <= 16'h0FAE;    16'd50498: out <= 16'h061A;    16'd50499: out <= 16'h06C1;
    16'd50500: out <= 16'h020B;    16'd50501: out <= 16'h03FB;    16'd50502: out <= 16'h05C0;    16'd50503: out <= 16'h02E4;
    16'd50504: out <= 16'hFEDC;    16'd50505: out <= 16'hFF90;    16'd50506: out <= 16'h02CC;    16'd50507: out <= 16'h032E;
    16'd50508: out <= 16'h0379;    16'd50509: out <= 16'h0413;    16'd50510: out <= 16'hFEB8;    16'd50511: out <= 16'h056D;
    16'd50512: out <= 16'h053F;    16'd50513: out <= 16'h0117;    16'd50514: out <= 16'h0155;    16'd50515: out <= 16'h0536;
    16'd50516: out <= 16'h0898;    16'd50517: out <= 16'h0B1C;    16'd50518: out <= 16'h0670;    16'd50519: out <= 16'h0138;
    16'd50520: out <= 16'h0339;    16'd50521: out <= 16'h0312;    16'd50522: out <= 16'hFF5F;    16'd50523: out <= 16'h03B8;
    16'd50524: out <= 16'h020B;    16'd50525: out <= 16'h03FF;    16'd50526: out <= 16'h0326;    16'd50527: out <= 16'hFFEF;
    16'd50528: out <= 16'h00C2;    16'd50529: out <= 16'h01AE;    16'd50530: out <= 16'h0517;    16'd50531: out <= 16'h000F;
    16'd50532: out <= 16'h0365;    16'd50533: out <= 16'h043C;    16'd50534: out <= 16'h0432;    16'd50535: out <= 16'h066C;
    16'd50536: out <= 16'h0664;    16'd50537: out <= 16'h06D8;    16'd50538: out <= 16'hFEF2;    16'd50539: out <= 16'hFDB8;
    16'd50540: out <= 16'hFB71;    16'd50541: out <= 16'h0C21;    16'd50542: out <= 16'hFC87;    16'd50543: out <= 16'h0650;
    16'd50544: out <= 16'h03D4;    16'd50545: out <= 16'h042B;    16'd50546: out <= 16'h0608;    16'd50547: out <= 16'hFC09;
    16'd50548: out <= 16'h06FF;    16'd50549: out <= 16'hFF66;    16'd50550: out <= 16'hFFC1;    16'd50551: out <= 16'h0581;
    16'd50552: out <= 16'h04D3;    16'd50553: out <= 16'hFBEB;    16'd50554: out <= 16'hFDF6;    16'd50555: out <= 16'h0346;
    16'd50556: out <= 16'h0092;    16'd50557: out <= 16'h05D4;    16'd50558: out <= 16'h0C1D;    16'd50559: out <= 16'hF940;
    16'd50560: out <= 16'h028C;    16'd50561: out <= 16'h0564;    16'd50562: out <= 16'h06E5;    16'd50563: out <= 16'hFFAA;
    16'd50564: out <= 16'h0D01;    16'd50565: out <= 16'h0698;    16'd50566: out <= 16'hFFB2;    16'd50567: out <= 16'h0476;
    16'd50568: out <= 16'h0704;    16'd50569: out <= 16'h0111;    16'd50570: out <= 16'h0715;    16'd50571: out <= 16'hFD63;
    16'd50572: out <= 16'h03A5;    16'd50573: out <= 16'h0029;    16'd50574: out <= 16'h0490;    16'd50575: out <= 16'h03B8;
    16'd50576: out <= 16'h0B7E;    16'd50577: out <= 16'hFEE5;    16'd50578: out <= 16'h002C;    16'd50579: out <= 16'hFF3B;
    16'd50580: out <= 16'h0172;    16'd50581: out <= 16'h00C0;    16'd50582: out <= 16'h0327;    16'd50583: out <= 16'h00CB;
    16'd50584: out <= 16'h02C4;    16'd50585: out <= 16'h05AE;    16'd50586: out <= 16'h0631;    16'd50587: out <= 16'h09C4;
    16'd50588: out <= 16'h0926;    16'd50589: out <= 16'hFDFB;    16'd50590: out <= 16'hFE08;    16'd50591: out <= 16'h0359;
    16'd50592: out <= 16'hFF17;    16'd50593: out <= 16'h036A;    16'd50594: out <= 16'h0714;    16'd50595: out <= 16'h021A;
    16'd50596: out <= 16'h01BF;    16'd50597: out <= 16'hF8FE;    16'd50598: out <= 16'h03D5;    16'd50599: out <= 16'h08E2;
    16'd50600: out <= 16'hFF95;    16'd50601: out <= 16'h0239;    16'd50602: out <= 16'h0145;    16'd50603: out <= 16'h0322;
    16'd50604: out <= 16'h06F9;    16'd50605: out <= 16'h0890;    16'd50606: out <= 16'h0398;    16'd50607: out <= 16'h02A2;
    16'd50608: out <= 16'h04AB;    16'd50609: out <= 16'h03BE;    16'd50610: out <= 16'h0786;    16'd50611: out <= 16'h07B4;
    16'd50612: out <= 16'h020F;    16'd50613: out <= 16'h0735;    16'd50614: out <= 16'h03BB;    16'd50615: out <= 16'h040E;
    16'd50616: out <= 16'h04F7;    16'd50617: out <= 16'hFD03;    16'd50618: out <= 16'h014C;    16'd50619: out <= 16'hFE8E;
    16'd50620: out <= 16'h019C;    16'd50621: out <= 16'h00ED;    16'd50622: out <= 16'h077D;    16'd50623: out <= 16'h058E;
    16'd50624: out <= 16'h0520;    16'd50625: out <= 16'h05D0;    16'd50626: out <= 16'hFFCA;    16'd50627: out <= 16'h0061;
    16'd50628: out <= 16'hFC26;    16'd50629: out <= 16'hFCA8;    16'd50630: out <= 16'h00B6;    16'd50631: out <= 16'h0077;
    16'd50632: out <= 16'h040E;    16'd50633: out <= 16'hFBF0;    16'd50634: out <= 16'h0229;    16'd50635: out <= 16'hFD64;
    16'd50636: out <= 16'hFB4A;    16'd50637: out <= 16'h0037;    16'd50638: out <= 16'h031D;    16'd50639: out <= 16'hFD63;
    16'd50640: out <= 16'hF7E5;    16'd50641: out <= 16'h011C;    16'd50642: out <= 16'h037F;    16'd50643: out <= 16'h0063;
    16'd50644: out <= 16'h0541;    16'd50645: out <= 16'hF80A;    16'd50646: out <= 16'hFF5B;    16'd50647: out <= 16'h01FB;
    16'd50648: out <= 16'h043B;    16'd50649: out <= 16'h007B;    16'd50650: out <= 16'hFE06;    16'd50651: out <= 16'hF9C7;
    16'd50652: out <= 16'hFD56;    16'd50653: out <= 16'hFED1;    16'd50654: out <= 16'h044B;    16'd50655: out <= 16'h0395;
    16'd50656: out <= 16'h0002;    16'd50657: out <= 16'hFDF3;    16'd50658: out <= 16'hFB3F;    16'd50659: out <= 16'hFEF5;
    16'd50660: out <= 16'h0319;    16'd50661: out <= 16'h051A;    16'd50662: out <= 16'h05A1;    16'd50663: out <= 16'h038F;
    16'd50664: out <= 16'h0361;    16'd50665: out <= 16'h0195;    16'd50666: out <= 16'h018C;    16'd50667: out <= 16'hFCBB;
    16'd50668: out <= 16'hFDBA;    16'd50669: out <= 16'hFB83;    16'd50670: out <= 16'h04BE;    16'd50671: out <= 16'h0092;
    16'd50672: out <= 16'h022E;    16'd50673: out <= 16'h0205;    16'd50674: out <= 16'h0287;    16'd50675: out <= 16'hFD24;
    16'd50676: out <= 16'hFA4F;    16'd50677: out <= 16'h02CB;    16'd50678: out <= 16'h0248;    16'd50679: out <= 16'h0070;
    16'd50680: out <= 16'hFF87;    16'd50681: out <= 16'h0141;    16'd50682: out <= 16'hFC28;    16'd50683: out <= 16'hFDF6;
    16'd50684: out <= 16'h0081;    16'd50685: out <= 16'h0121;    16'd50686: out <= 16'hFEDB;    16'd50687: out <= 16'h02D7;
    16'd50688: out <= 16'hFD8C;    16'd50689: out <= 16'h0232;    16'd50690: out <= 16'h05BB;    16'd50691: out <= 16'h01E4;
    16'd50692: out <= 16'hF853;    16'd50693: out <= 16'hFF26;    16'd50694: out <= 16'hFFD8;    16'd50695: out <= 16'h0271;
    16'd50696: out <= 16'hFDB6;    16'd50697: out <= 16'hF8DE;    16'd50698: out <= 16'hFCC3;    16'd50699: out <= 16'hFF10;
    16'd50700: out <= 16'hFC6D;    16'd50701: out <= 16'h0585;    16'd50702: out <= 16'hFACB;    16'd50703: out <= 16'h024E;
    16'd50704: out <= 16'h0153;    16'd50705: out <= 16'h03AC;    16'd50706: out <= 16'hFECF;    16'd50707: out <= 16'h0271;
    16'd50708: out <= 16'h02AD;    16'd50709: out <= 16'h0123;    16'd50710: out <= 16'h0778;    16'd50711: out <= 16'h00BA;
    16'd50712: out <= 16'hFD3C;    16'd50713: out <= 16'h05DD;    16'd50714: out <= 16'h02F6;    16'd50715: out <= 16'h00E0;
    16'd50716: out <= 16'hFB3F;    16'd50717: out <= 16'h00AB;    16'd50718: out <= 16'h01F4;    16'd50719: out <= 16'hFA2F;
    16'd50720: out <= 16'h045A;    16'd50721: out <= 16'hFEA7;    16'd50722: out <= 16'h080E;    16'd50723: out <= 16'hFAEA;
    16'd50724: out <= 16'h0514;    16'd50725: out <= 16'h038E;    16'd50726: out <= 16'h035C;    16'd50727: out <= 16'h0362;
    16'd50728: out <= 16'h0143;    16'd50729: out <= 16'hFADD;    16'd50730: out <= 16'h0056;    16'd50731: out <= 16'h03B7;
    16'd50732: out <= 16'h0387;    16'd50733: out <= 16'h02F8;    16'd50734: out <= 16'h047A;    16'd50735: out <= 16'h056D;
    16'd50736: out <= 16'hFD97;    16'd50737: out <= 16'h0429;    16'd50738: out <= 16'h070F;    16'd50739: out <= 16'h01AB;
    16'd50740: out <= 16'h07BA;    16'd50741: out <= 16'h07EC;    16'd50742: out <= 16'h055D;    16'd50743: out <= 16'h02B2;
    16'd50744: out <= 16'hF99B;    16'd50745: out <= 16'hFE6C;    16'd50746: out <= 16'h0838;    16'd50747: out <= 16'h0143;
    16'd50748: out <= 16'h06B7;    16'd50749: out <= 16'h0066;    16'd50750: out <= 16'hFE13;    16'd50751: out <= 16'h0685;
    16'd50752: out <= 16'h0374;    16'd50753: out <= 16'h0527;    16'd50754: out <= 16'h0706;    16'd50755: out <= 16'hFECA;
    16'd50756: out <= 16'h02C7;    16'd50757: out <= 16'h001A;    16'd50758: out <= 16'hF9F8;    16'd50759: out <= 16'h0135;
    16'd50760: out <= 16'h0A86;    16'd50761: out <= 16'h05FF;    16'd50762: out <= 16'h04D1;    16'd50763: out <= 16'h0904;
    16'd50764: out <= 16'h0051;    16'd50765: out <= 16'h018B;    16'd50766: out <= 16'h04EA;    16'd50767: out <= 16'h0807;
    16'd50768: out <= 16'h00E6;    16'd50769: out <= 16'hFF95;    16'd50770: out <= 16'h081C;    16'd50771: out <= 16'h061D;
    16'd50772: out <= 16'h04A6;    16'd50773: out <= 16'h00E3;    16'd50774: out <= 16'hFFBA;    16'd50775: out <= 16'h0659;
    16'd50776: out <= 16'h0AAE;    16'd50777: out <= 16'h0A2C;    16'd50778: out <= 16'h08F5;    16'd50779: out <= 16'h004F;
    16'd50780: out <= 16'h03B7;    16'd50781: out <= 16'h0565;    16'd50782: out <= 16'h089C;    16'd50783: out <= 16'h09E3;
    16'd50784: out <= 16'h0400;    16'd50785: out <= 16'h03CC;    16'd50786: out <= 16'h080B;    16'd50787: out <= 16'h0271;
    16'd50788: out <= 16'hFF98;    16'd50789: out <= 16'h061B;    16'd50790: out <= 16'h01CB;    16'd50791: out <= 16'hFFBB;
    16'd50792: out <= 16'hFBDA;    16'd50793: out <= 16'hFC39;    16'd50794: out <= 16'h02CF;    16'd50795: out <= 16'hFA29;
    16'd50796: out <= 16'h0017;    16'd50797: out <= 16'h013B;    16'd50798: out <= 16'h017C;    16'd50799: out <= 16'hFF0A;
    16'd50800: out <= 16'h03CC;    16'd50801: out <= 16'h023D;    16'd50802: out <= 16'h097F;    16'd50803: out <= 16'h04FA;
    16'd50804: out <= 16'hFCFF;    16'd50805: out <= 16'h0006;    16'd50806: out <= 16'h03B7;    16'd50807: out <= 16'h0044;
    16'd50808: out <= 16'hF81D;    16'd50809: out <= 16'hFD4A;    16'd50810: out <= 16'h07FC;    16'd50811: out <= 16'hFC11;
    16'd50812: out <= 16'h035F;    16'd50813: out <= 16'h002A;    16'd50814: out <= 16'hFEB4;    16'd50815: out <= 16'h006E;
    16'd50816: out <= 16'h047D;    16'd50817: out <= 16'h0901;    16'd50818: out <= 16'h053A;    16'd50819: out <= 16'h0768;
    16'd50820: out <= 16'hFBE7;    16'd50821: out <= 16'h02D1;    16'd50822: out <= 16'h0304;    16'd50823: out <= 16'hFCE9;
    16'd50824: out <= 16'h0324;    16'd50825: out <= 16'hFA68;    16'd50826: out <= 16'h0791;    16'd50827: out <= 16'h07BF;
    16'd50828: out <= 16'h06B7;    16'd50829: out <= 16'h020B;    16'd50830: out <= 16'h0588;    16'd50831: out <= 16'h0965;
    16'd50832: out <= 16'h073A;    16'd50833: out <= 16'h0226;    16'd50834: out <= 16'h07A2;    16'd50835: out <= 16'h0621;
    16'd50836: out <= 16'hFDBA;    16'd50837: out <= 16'hFCAB;    16'd50838: out <= 16'hFCB8;    16'd50839: out <= 16'h03B4;
    16'd50840: out <= 16'h05BD;    16'd50841: out <= 16'hFED2;    16'd50842: out <= 16'h00E6;    16'd50843: out <= 16'h0296;
    16'd50844: out <= 16'h053B;    16'd50845: out <= 16'hFFC8;    16'd50846: out <= 16'h03E7;    16'd50847: out <= 16'h0618;
    16'd50848: out <= 16'h03F4;    16'd50849: out <= 16'h0203;    16'd50850: out <= 16'h06A2;    16'd50851: out <= 16'h06C2;
    16'd50852: out <= 16'h05E8;    16'd50853: out <= 16'h06FD;    16'd50854: out <= 16'h076C;    16'd50855: out <= 16'h026C;
    16'd50856: out <= 16'h061A;    16'd50857: out <= 16'h03BF;    16'd50858: out <= 16'h083E;    16'd50859: out <= 16'h02C4;
    16'd50860: out <= 16'hFF51;    16'd50861: out <= 16'h0138;    16'd50862: out <= 16'h0147;    16'd50863: out <= 16'h05BC;
    16'd50864: out <= 16'h03B8;    16'd50865: out <= 16'h0066;    16'd50866: out <= 16'h03C8;    16'd50867: out <= 16'h02F9;
    16'd50868: out <= 16'h02B1;    16'd50869: out <= 16'h08DE;    16'd50870: out <= 16'hFDF4;    16'd50871: out <= 16'hFD9C;
    16'd50872: out <= 16'h05D7;    16'd50873: out <= 16'h00D3;    16'd50874: out <= 16'h02BD;    16'd50875: out <= 16'h02DB;
    16'd50876: out <= 16'hFF03;    16'd50877: out <= 16'h0799;    16'd50878: out <= 16'h043C;    16'd50879: out <= 16'h02B1;
    16'd50880: out <= 16'h01F6;    16'd50881: out <= 16'h039C;    16'd50882: out <= 16'h013D;    16'd50883: out <= 16'h0115;
    16'd50884: out <= 16'hFFA2;    16'd50885: out <= 16'hF8B0;    16'd50886: out <= 16'hFACD;    16'd50887: out <= 16'hFD5A;
    16'd50888: out <= 16'hFFAD;    16'd50889: out <= 16'hFE0C;    16'd50890: out <= 16'h0107;    16'd50891: out <= 16'h0CE0;
    16'd50892: out <= 16'h0045;    16'd50893: out <= 16'h03A4;    16'd50894: out <= 16'hFF07;    16'd50895: out <= 16'hF8AF;
    16'd50896: out <= 16'hFE70;    16'd50897: out <= 16'hFEB3;    16'd50898: out <= 16'h07E0;    16'd50899: out <= 16'hFF52;
    16'd50900: out <= 16'h046E;    16'd50901: out <= 16'hFFFB;    16'd50902: out <= 16'h053B;    16'd50903: out <= 16'h0233;
    16'd50904: out <= 16'hFF87;    16'd50905: out <= 16'h06EB;    16'd50906: out <= 16'hFF4D;    16'd50907: out <= 16'h0168;
    16'd50908: out <= 16'h01DC;    16'd50909: out <= 16'h0462;    16'd50910: out <= 16'h00BC;    16'd50911: out <= 16'hFBBE;
    16'd50912: out <= 16'h0335;    16'd50913: out <= 16'hFF0C;    16'd50914: out <= 16'hFEE4;    16'd50915: out <= 16'hFB7A;
    16'd50916: out <= 16'hFA44;    16'd50917: out <= 16'hFD83;    16'd50918: out <= 16'hFF90;    16'd50919: out <= 16'hFEE7;
    16'd50920: out <= 16'h053C;    16'd50921: out <= 16'h0315;    16'd50922: out <= 16'h0222;    16'd50923: out <= 16'h054B;
    16'd50924: out <= 16'hFD3D;    16'd50925: out <= 16'hFBB7;    16'd50926: out <= 16'hFAF5;    16'd50927: out <= 16'hFE08;
    16'd50928: out <= 16'hF73E;    16'd50929: out <= 16'h02D7;    16'd50930: out <= 16'hFFA0;    16'd50931: out <= 16'hFB5B;
    16'd50932: out <= 16'hFB5A;    16'd50933: out <= 16'h034B;    16'd50934: out <= 16'hF994;    16'd50935: out <= 16'hFCAB;
    16'd50936: out <= 16'hFC4A;    16'd50937: out <= 16'h0249;    16'd50938: out <= 16'h0433;    16'd50939: out <= 16'hFC94;
    16'd50940: out <= 16'h018B;    16'd50941: out <= 16'h06CE;    16'd50942: out <= 16'hFCB7;    16'd50943: out <= 16'h0141;
    16'd50944: out <= 16'hF4C8;    16'd50945: out <= 16'h025E;    16'd50946: out <= 16'hFD28;    16'd50947: out <= 16'hFE77;
    16'd50948: out <= 16'hFEBE;    16'd50949: out <= 16'hFC4C;    16'd50950: out <= 16'hF867;    16'd50951: out <= 16'h01D1;
    16'd50952: out <= 16'hFD80;    16'd50953: out <= 16'hFD29;    16'd50954: out <= 16'hFE42;    16'd50955: out <= 16'hFC96;
    16'd50956: out <= 16'hFAA3;    16'd50957: out <= 16'hFFFA;    16'd50958: out <= 16'hFC53;    16'd50959: out <= 16'h02B9;
    16'd50960: out <= 16'h04BD;    16'd50961: out <= 16'hFF94;    16'd50962: out <= 16'h045A;    16'd50963: out <= 16'h027B;
    16'd50964: out <= 16'hFED5;    16'd50965: out <= 16'hFF16;    16'd50966: out <= 16'h02B1;    16'd50967: out <= 16'hFB73;
    16'd50968: out <= 16'hFA38;    16'd50969: out <= 16'hFA76;    16'd50970: out <= 16'hFE6E;    16'd50971: out <= 16'h0163;
    16'd50972: out <= 16'hFF16;    16'd50973: out <= 16'h02F5;    16'd50974: out <= 16'h058B;    16'd50975: out <= 16'hF948;
    16'd50976: out <= 16'h0038;    16'd50977: out <= 16'hFDD0;    16'd50978: out <= 16'h0647;    16'd50979: out <= 16'h0384;
    16'd50980: out <= 16'h01E6;    16'd50981: out <= 16'h0013;    16'd50982: out <= 16'h0421;    16'd50983: out <= 16'h00AB;
    16'd50984: out <= 16'h0158;    16'd50985: out <= 16'h00A8;    16'd50986: out <= 16'h0385;    16'd50987: out <= 16'h00DC;
    16'd50988: out <= 16'h079A;    16'd50989: out <= 16'hFD3A;    16'd50990: out <= 16'h0C92;    16'd50991: out <= 16'h07F0;
    16'd50992: out <= 16'h04AA;    16'd50993: out <= 16'h0CE2;    16'd50994: out <= 16'h023C;    16'd50995: out <= 16'h076A;
    16'd50996: out <= 16'h061F;    16'd50997: out <= 16'h06A3;    16'd50998: out <= 16'h0658;    16'd50999: out <= 16'h0945;
    16'd51000: out <= 16'h0115;    16'd51001: out <= 16'h0588;    16'd51002: out <= 16'hFD11;    16'd51003: out <= 16'h0AB9;
    16'd51004: out <= 16'h024A;    16'd51005: out <= 16'h0081;    16'd51006: out <= 16'h02F2;    16'd51007: out <= 16'h06C6;
    16'd51008: out <= 16'h04F0;    16'd51009: out <= 16'h03F1;    16'd51010: out <= 16'h0AEC;    16'd51011: out <= 16'h0571;
    16'd51012: out <= 16'h00DE;    16'd51013: out <= 16'h07E9;    16'd51014: out <= 16'h0641;    16'd51015: out <= 16'h0181;
    16'd51016: out <= 16'h069B;    16'd51017: out <= 16'h0508;    16'd51018: out <= 16'h0533;    16'd51019: out <= 16'h00F2;
    16'd51020: out <= 16'h04A6;    16'd51021: out <= 16'h002A;    16'd51022: out <= 16'h0285;    16'd51023: out <= 16'h0281;
    16'd51024: out <= 16'h0576;    16'd51025: out <= 16'h027E;    16'd51026: out <= 16'h0651;    16'd51027: out <= 16'h0650;
    16'd51028: out <= 16'h0835;    16'd51029: out <= 16'h08D4;    16'd51030: out <= 16'h06BC;    16'd51031: out <= 16'h0414;
    16'd51032: out <= 16'hFD09;    16'd51033: out <= 16'h04A4;    16'd51034: out <= 16'h0114;    16'd51035: out <= 16'h086D;
    16'd51036: out <= 16'h0750;    16'd51037: out <= 16'h038A;    16'd51038: out <= 16'h090B;    16'd51039: out <= 16'h0485;
    16'd51040: out <= 16'h055D;    16'd51041: out <= 16'h0066;    16'd51042: out <= 16'h0215;    16'd51043: out <= 16'h028F;
    16'd51044: out <= 16'h0821;    16'd51045: out <= 16'hFE99;    16'd51046: out <= 16'hFECA;    16'd51047: out <= 16'h085B;
    16'd51048: out <= 16'h0847;    16'd51049: out <= 16'h0715;    16'd51050: out <= 16'hFD2C;    16'd51051: out <= 16'hFEA1;
    16'd51052: out <= 16'h04D9;    16'd51053: out <= 16'h01A2;    16'd51054: out <= 16'hFF6E;    16'd51055: out <= 16'h00A2;
    16'd51056: out <= 16'h01D1;    16'd51057: out <= 16'h001F;    16'd51058: out <= 16'h01C4;    16'd51059: out <= 16'hFC16;
    16'd51060: out <= 16'hF841;    16'd51061: out <= 16'hFACD;    16'd51062: out <= 16'hFB90;    16'd51063: out <= 16'hFF0A;
    16'd51064: out <= 16'h0387;    16'd51065: out <= 16'h0122;    16'd51066: out <= 16'hFEFA;    16'd51067: out <= 16'h04A7;
    16'd51068: out <= 16'h0195;    16'd51069: out <= 16'h01DF;    16'd51070: out <= 16'h04BC;    16'd51071: out <= 16'h02B8;
    16'd51072: out <= 16'hFCD5;    16'd51073: out <= 16'h0761;    16'd51074: out <= 16'h09BF;    16'd51075: out <= 16'h074B;
    16'd51076: out <= 16'h030F;    16'd51077: out <= 16'h08A3;    16'd51078: out <= 16'h033D;    16'd51079: out <= 16'h0984;
    16'd51080: out <= 16'h0BFC;    16'd51081: out <= 16'h0BD9;    16'd51082: out <= 16'h005D;    16'd51083: out <= 16'h09C1;
    16'd51084: out <= 16'h089C;    16'd51085: out <= 16'h0234;    16'd51086: out <= 16'h03BD;    16'd51087: out <= 16'h072C;
    16'd51088: out <= 16'h03FC;    16'd51089: out <= 16'h04F0;    16'd51090: out <= 16'h0508;    16'd51091: out <= 16'h067A;
    16'd51092: out <= 16'h055C;    16'd51093: out <= 16'hFC20;    16'd51094: out <= 16'h051B;    16'd51095: out <= 16'hF8F8;
    16'd51096: out <= 16'h0B4F;    16'd51097: out <= 16'h0393;    16'd51098: out <= 16'h01C3;    16'd51099: out <= 16'hFF0D;
    16'd51100: out <= 16'h0621;    16'd51101: out <= 16'h03D3;    16'd51102: out <= 16'h0208;    16'd51103: out <= 16'h07B3;
    16'd51104: out <= 16'h0948;    16'd51105: out <= 16'h0230;    16'd51106: out <= 16'h00ED;    16'd51107: out <= 16'h025A;
    16'd51108: out <= 16'h06C9;    16'd51109: out <= 16'h0728;    16'd51110: out <= 16'h08E4;    16'd51111: out <= 16'h055F;
    16'd51112: out <= 16'h04D1;    16'd51113: out <= 16'h029E;    16'd51114: out <= 16'h0431;    16'd51115: out <= 16'h04BA;
    16'd51116: out <= 16'h00CE;    16'd51117: out <= 16'hFFA9;    16'd51118: out <= 16'h03B7;    16'd51119: out <= 16'h008B;
    16'd51120: out <= 16'h027F;    16'd51121: out <= 16'hFDF3;    16'd51122: out <= 16'h0861;    16'd51123: out <= 16'h03ED;
    16'd51124: out <= 16'h054F;    16'd51125: out <= 16'h0687;    16'd51126: out <= 16'h02E8;    16'd51127: out <= 16'h017C;
    16'd51128: out <= 16'h0199;    16'd51129: out <= 16'h094F;    16'd51130: out <= 16'h00A3;    16'd51131: out <= 16'h02A9;
    16'd51132: out <= 16'h0547;    16'd51133: out <= 16'h0169;    16'd51134: out <= 16'h0224;    16'd51135: out <= 16'h013A;
    16'd51136: out <= 16'hFA47;    16'd51137: out <= 16'h0175;    16'd51138: out <= 16'h05FF;    16'd51139: out <= 16'h06B0;
    16'd51140: out <= 16'hFBEB;    16'd51141: out <= 16'hFFAB;    16'd51142: out <= 16'hFFF7;    16'd51143: out <= 16'h042C;
    16'd51144: out <= 16'h01E2;    16'd51145: out <= 16'hFC48;    16'd51146: out <= 16'h04D4;    16'd51147: out <= 16'h0250;
    16'd51148: out <= 16'h06A1;    16'd51149: out <= 16'h03FD;    16'd51150: out <= 16'hF997;    16'd51151: out <= 16'h04D0;
    16'd51152: out <= 16'h06A8;    16'd51153: out <= 16'h06E2;    16'd51154: out <= 16'h08A8;    16'd51155: out <= 16'hFC83;
    16'd51156: out <= 16'hFF14;    16'd51157: out <= 16'hFF75;    16'd51158: out <= 16'hFD26;    16'd51159: out <= 16'hF988;
    16'd51160: out <= 16'hFF2F;    16'd51161: out <= 16'h0106;    16'd51162: out <= 16'hFCB9;    16'd51163: out <= 16'hFF33;
    16'd51164: out <= 16'hFB9E;    16'd51165: out <= 16'h03CB;    16'd51166: out <= 16'h038F;    16'd51167: out <= 16'hF417;
    16'd51168: out <= 16'h0111;    16'd51169: out <= 16'hFF93;    16'd51170: out <= 16'h02CB;    16'd51171: out <= 16'h07EB;
    16'd51172: out <= 16'h0251;    16'd51173: out <= 16'h0593;    16'd51174: out <= 16'hFE6B;    16'd51175: out <= 16'hFF18;
    16'd51176: out <= 16'hF9E1;    16'd51177: out <= 16'h02F6;    16'd51178: out <= 16'hFEC2;    16'd51179: out <= 16'hF87A;
    16'd51180: out <= 16'h03BE;    16'd51181: out <= 16'h0AE1;    16'd51182: out <= 16'h0549;    16'd51183: out <= 16'hFF28;
    16'd51184: out <= 16'hFB9E;    16'd51185: out <= 16'h02D9;    16'd51186: out <= 16'hFFD8;    16'd51187: out <= 16'h033E;
    16'd51188: out <= 16'h0228;    16'd51189: out <= 16'h0399;    16'd51190: out <= 16'hFB0F;    16'd51191: out <= 16'h00C1;
    16'd51192: out <= 16'hFC6B;    16'd51193: out <= 16'hFF94;    16'd51194: out <= 16'h037B;    16'd51195: out <= 16'hFF27;
    16'd51196: out <= 16'h0422;    16'd51197: out <= 16'hFEE0;    16'd51198: out <= 16'hFF45;    16'd51199: out <= 16'h01D9;
    16'd51200: out <= 16'hFD74;    16'd51201: out <= 16'h0034;    16'd51202: out <= 16'hFE69;    16'd51203: out <= 16'h008D;
    16'd51204: out <= 16'h02F0;    16'd51205: out <= 16'hF90A;    16'd51206: out <= 16'h0645;    16'd51207: out <= 16'hF806;
    16'd51208: out <= 16'hFBFE;    16'd51209: out <= 16'h02E2;    16'd51210: out <= 16'h0258;    16'd51211: out <= 16'h0292;
    16'd51212: out <= 16'h0173;    16'd51213: out <= 16'hFBAA;    16'd51214: out <= 16'h02A4;    16'd51215: out <= 16'h0593;
    16'd51216: out <= 16'h01E9;    16'd51217: out <= 16'h00A4;    16'd51218: out <= 16'h0459;    16'd51219: out <= 16'hFB0D;
    16'd51220: out <= 16'h0694;    16'd51221: out <= 16'h0A70;    16'd51222: out <= 16'h0196;    16'd51223: out <= 16'hFEE9;
    16'd51224: out <= 16'hF8BC;    16'd51225: out <= 16'hFD82;    16'd51226: out <= 16'hFDC6;    16'd51227: out <= 16'h02CE;
    16'd51228: out <= 16'h00E5;    16'd51229: out <= 16'hFE66;    16'd51230: out <= 16'hF4EB;    16'd51231: out <= 16'hFB13;
    16'd51232: out <= 16'h0273;    16'd51233: out <= 16'h024C;    16'd51234: out <= 16'h0067;    16'd51235: out <= 16'hFE00;
    16'd51236: out <= 16'h0090;    16'd51237: out <= 16'h0287;    16'd51238: out <= 16'h00D0;    16'd51239: out <= 16'hFFE0;
    16'd51240: out <= 16'hFC71;    16'd51241: out <= 16'hFFF5;    16'd51242: out <= 16'h0397;    16'd51243: out <= 16'hFEBD;
    16'd51244: out <= 16'h05FA;    16'd51245: out <= 16'h0375;    16'd51246: out <= 16'h063E;    16'd51247: out <= 16'h040D;
    16'd51248: out <= 16'hFF85;    16'd51249: out <= 16'h003D;    16'd51250: out <= 16'h0882;    16'd51251: out <= 16'h04F4;
    16'd51252: out <= 16'h0027;    16'd51253: out <= 16'hFED2;    16'd51254: out <= 16'h04E3;    16'd51255: out <= 16'hFB06;
    16'd51256: out <= 16'h0231;    16'd51257: out <= 16'h05DF;    16'd51258: out <= 16'h052C;    16'd51259: out <= 16'h0A95;
    16'd51260: out <= 16'hFF30;    16'd51261: out <= 16'h0206;    16'd51262: out <= 16'h04F9;    16'd51263: out <= 16'h05B0;
    16'd51264: out <= 16'h0497;    16'd51265: out <= 16'hFF7F;    16'd51266: out <= 16'h029B;    16'd51267: out <= 16'h0268;
    16'd51268: out <= 16'h006B;    16'd51269: out <= 16'h050E;    16'd51270: out <= 16'h0489;    16'd51271: out <= 16'h008B;
    16'd51272: out <= 16'h0087;    16'd51273: out <= 16'hFF59;    16'd51274: out <= 16'hFFF3;    16'd51275: out <= 16'h03D5;
    16'd51276: out <= 16'h00E4;    16'd51277: out <= 16'h03CC;    16'd51278: out <= 16'h02C1;    16'd51279: out <= 16'hFFA4;
    16'd51280: out <= 16'h09E5;    16'd51281: out <= 16'h0A98;    16'd51282: out <= 16'h0989;    16'd51283: out <= 16'h00D4;
    16'd51284: out <= 16'h04F4;    16'd51285: out <= 16'hFB64;    16'd51286: out <= 16'h044B;    16'd51287: out <= 16'h06DB;
    16'd51288: out <= 16'h00C7;    16'd51289: out <= 16'h0373;    16'd51290: out <= 16'h0297;    16'd51291: out <= 16'hFF0F;
    16'd51292: out <= 16'hFE4F;    16'd51293: out <= 16'hFEC9;    16'd51294: out <= 16'h05E3;    16'd51295: out <= 16'hFF8E;
    16'd51296: out <= 16'hFEE7;    16'd51297: out <= 16'h0709;    16'd51298: out <= 16'h03E5;    16'd51299: out <= 16'h0880;
    16'd51300: out <= 16'h0204;    16'd51301: out <= 16'h0455;    16'd51302: out <= 16'h042C;    16'd51303: out <= 16'h018E;
    16'd51304: out <= 16'h0213;    16'd51305: out <= 16'h0366;    16'd51306: out <= 16'hFF61;    16'd51307: out <= 16'hFE92;
    16'd51308: out <= 16'hFEF3;    16'd51309: out <= 16'hFE93;    16'd51310: out <= 16'h045D;    16'd51311: out <= 16'h00FF;
    16'd51312: out <= 16'hFEF5;    16'd51313: out <= 16'h018C;    16'd51314: out <= 16'hFD9F;    16'd51315: out <= 16'hFCCD;
    16'd51316: out <= 16'hFE67;    16'd51317: out <= 16'hFD85;    16'd51318: out <= 16'hFDCC;    16'd51319: out <= 16'hFEC8;
    16'd51320: out <= 16'h00A2;    16'd51321: out <= 16'h0986;    16'd51322: out <= 16'hFC60;    16'd51323: out <= 16'hFE37;
    16'd51324: out <= 16'h05C8;    16'd51325: out <= 16'h0729;    16'd51326: out <= 16'h0596;    16'd51327: out <= 16'h03F8;
    16'd51328: out <= 16'h09A8;    16'd51329: out <= 16'h0298;    16'd51330: out <= 16'hFEC0;    16'd51331: out <= 16'h0313;
    16'd51332: out <= 16'h0389;    16'd51333: out <= 16'h06EF;    16'd51334: out <= 16'h07E7;    16'd51335: out <= 16'h01E6;
    16'd51336: out <= 16'h0111;    16'd51337: out <= 16'h0328;    16'd51338: out <= 16'h0945;    16'd51339: out <= 16'h0A1F;
    16'd51340: out <= 16'h0634;    16'd51341: out <= 16'hFE60;    16'd51342: out <= 16'h032D;    16'd51343: out <= 16'h026E;
    16'd51344: out <= 16'h044A;    16'd51345: out <= 16'h0587;    16'd51346: out <= 16'h0759;    16'd51347: out <= 16'h04AE;
    16'd51348: out <= 16'h0528;    16'd51349: out <= 16'hFE68;    16'd51350: out <= 16'h00E1;    16'd51351: out <= 16'h0A66;
    16'd51352: out <= 16'h027E;    16'd51353: out <= 16'h037C;    16'd51354: out <= 16'h08E8;    16'd51355: out <= 16'h0783;
    16'd51356: out <= 16'hFCC0;    16'd51357: out <= 16'h0690;    16'd51358: out <= 16'h01E9;    16'd51359: out <= 16'h0476;
    16'd51360: out <= 16'hFFCE;    16'd51361: out <= 16'h0927;    16'd51362: out <= 16'h0627;    16'd51363: out <= 16'h0662;
    16'd51364: out <= 16'h0498;    16'd51365: out <= 16'h03F2;    16'd51366: out <= 16'h01F5;    16'd51367: out <= 16'h04B8;
    16'd51368: out <= 16'h02D2;    16'd51369: out <= 16'h07C6;    16'd51370: out <= 16'h01EE;    16'd51371: out <= 16'h039D;
    16'd51372: out <= 16'h071F;    16'd51373: out <= 16'h0473;    16'd51374: out <= 16'h0AA5;    16'd51375: out <= 16'h0455;
    16'd51376: out <= 16'h01B8;    16'd51377: out <= 16'h0458;    16'd51378: out <= 16'hFFA3;    16'd51379: out <= 16'h07EC;
    16'd51380: out <= 16'h026B;    16'd51381: out <= 16'h064D;    16'd51382: out <= 16'h0581;    16'd51383: out <= 16'h05FB;
    16'd51384: out <= 16'h05F4;    16'd51385: out <= 16'hFED1;    16'd51386: out <= 16'h033C;    16'd51387: out <= 16'hFBB6;
    16'd51388: out <= 16'h0344;    16'd51389: out <= 16'h0105;    16'd51390: out <= 16'h0417;    16'd51391: out <= 16'h081B;
    16'd51392: out <= 16'h06B5;    16'd51393: out <= 16'hFB1A;    16'd51394: out <= 16'hFFF4;    16'd51395: out <= 16'h0041;
    16'd51396: out <= 16'h0714;    16'd51397: out <= 16'hFCA9;    16'd51398: out <= 16'hFCC8;    16'd51399: out <= 16'hFE21;
    16'd51400: out <= 16'hFE1A;    16'd51401: out <= 16'hFF45;    16'd51402: out <= 16'h071A;    16'd51403: out <= 16'h0470;
    16'd51404: out <= 16'hFE83;    16'd51405: out <= 16'hFF95;    16'd51406: out <= 16'hFE3B;    16'd51407: out <= 16'h0221;
    16'd51408: out <= 16'hFEFD;    16'd51409: out <= 16'h026D;    16'd51410: out <= 16'hFE4C;    16'd51411: out <= 16'h058A;
    16'd51412: out <= 16'hFC08;    16'd51413: out <= 16'h05BF;    16'd51414: out <= 16'h05EE;    16'd51415: out <= 16'h03A9;
    16'd51416: out <= 16'hFC02;    16'd51417: out <= 16'h029A;    16'd51418: out <= 16'hFBD8;    16'd51419: out <= 16'h0201;
    16'd51420: out <= 16'h00FF;    16'd51421: out <= 16'h023F;    16'd51422: out <= 16'h0422;    16'd51423: out <= 16'hF98A;
    16'd51424: out <= 16'h02AB;    16'd51425: out <= 16'hFCC0;    16'd51426: out <= 16'hFB9B;    16'd51427: out <= 16'hFFB8;
    16'd51428: out <= 16'h011C;    16'd51429: out <= 16'hFCAF;    16'd51430: out <= 16'hFC02;    16'd51431: out <= 16'h0056;
    16'd51432: out <= 16'hFAB6;    16'd51433: out <= 16'hFA8D;    16'd51434: out <= 16'hFCEA;    16'd51435: out <= 16'hFE8D;
    16'd51436: out <= 16'h019B;    16'd51437: out <= 16'h0202;    16'd51438: out <= 16'hFC16;    16'd51439: out <= 16'h019C;
    16'd51440: out <= 16'h04DD;    16'd51441: out <= 16'hFDFF;    16'd51442: out <= 16'hFB41;    16'd51443: out <= 16'h0324;
    16'd51444: out <= 16'h05E0;    16'd51445: out <= 16'h0848;    16'd51446: out <= 16'h088F;    16'd51447: out <= 16'hFB88;
    16'd51448: out <= 16'hFF35;    16'd51449: out <= 16'hFDD6;    16'd51450: out <= 16'hFED1;    16'd51451: out <= 16'hF997;
    16'd51452: out <= 16'h0245;    16'd51453: out <= 16'hFD5F;    16'd51454: out <= 16'h00E0;    16'd51455: out <= 16'h033A;
    16'd51456: out <= 16'hFE7F;    16'd51457: out <= 16'hFCC3;    16'd51458: out <= 16'hFA00;    16'd51459: out <= 16'h01D0;
    16'd51460: out <= 16'h0243;    16'd51461: out <= 16'h09DE;    16'd51462: out <= 16'hFD80;    16'd51463: out <= 16'h051A;
    16'd51464: out <= 16'h0169;    16'd51465: out <= 16'hFA6D;    16'd51466: out <= 16'hFCDD;    16'd51467: out <= 16'hFA30;
    16'd51468: out <= 16'h00EE;    16'd51469: out <= 16'hFF86;    16'd51470: out <= 16'h03B0;    16'd51471: out <= 16'h0681;
    16'd51472: out <= 16'h01E1;    16'd51473: out <= 16'hFE44;    16'd51474: out <= 16'hFC0D;    16'd51475: out <= 16'hFFEE;
    16'd51476: out <= 16'hF7A1;    16'd51477: out <= 16'hFF69;    16'd51478: out <= 16'hFD90;    16'd51479: out <= 16'hF819;
    16'd51480: out <= 16'h038E;    16'd51481: out <= 16'hFD4C;    16'd51482: out <= 16'hFE78;    16'd51483: out <= 16'hFEFC;
    16'd51484: out <= 16'hFF4F;    16'd51485: out <= 16'hFF12;    16'd51486: out <= 16'h01F8;    16'd51487: out <= 16'h0301;
    16'd51488: out <= 16'h011B;    16'd51489: out <= 16'hFE92;    16'd51490: out <= 16'h00CD;    16'd51491: out <= 16'h010B;
    16'd51492: out <= 16'hFFBA;    16'd51493: out <= 16'h0140;    16'd51494: out <= 16'hFB5A;    16'd51495: out <= 16'h04D4;
    16'd51496: out <= 16'hFFA0;    16'd51497: out <= 16'hFD1E;    16'd51498: out <= 16'hFE6A;    16'd51499: out <= 16'hFF96;
    16'd51500: out <= 16'h034A;    16'd51501: out <= 16'h0441;    16'd51502: out <= 16'h0804;    16'd51503: out <= 16'hFB5C;
    16'd51504: out <= 16'h046D;    16'd51505: out <= 16'h0998;    16'd51506: out <= 16'hFF51;    16'd51507: out <= 16'h06D2;
    16'd51508: out <= 16'h02AF;    16'd51509: out <= 16'hFFE2;    16'd51510: out <= 16'h0DF0;    16'd51511: out <= 16'h08A5;
    16'd51512: out <= 16'hFDF5;    16'd51513: out <= 16'h0175;    16'd51514: out <= 16'h0888;    16'd51515: out <= 16'h0BB6;
    16'd51516: out <= 16'h0272;    16'd51517: out <= 16'hFF41;    16'd51518: out <= 16'h018E;    16'd51519: out <= 16'h0D94;
    16'd51520: out <= 16'h002A;    16'd51521: out <= 16'h01C0;    16'd51522: out <= 16'h0336;    16'd51523: out <= 16'h0A3E;
    16'd51524: out <= 16'h05F7;    16'd51525: out <= 16'h05B8;    16'd51526: out <= 16'h07FB;    16'd51527: out <= 16'h0513;
    16'd51528: out <= 16'h064B;    16'd51529: out <= 16'h0682;    16'd51530: out <= 16'h09BE;    16'd51531: out <= 16'h00EF;
    16'd51532: out <= 16'h08DA;    16'd51533: out <= 16'h0558;    16'd51534: out <= 16'h053A;    16'd51535: out <= 16'hFD5F;
    16'd51536: out <= 16'h0CAF;    16'd51537: out <= 16'h01D7;    16'd51538: out <= 16'h05FE;    16'd51539: out <= 16'h04B8;
    16'd51540: out <= 16'h050D;    16'd51541: out <= 16'hFFD6;    16'd51542: out <= 16'h0A65;    16'd51543: out <= 16'h039B;
    16'd51544: out <= 16'h09BD;    16'd51545: out <= 16'hFFF9;    16'd51546: out <= 16'hFD9B;    16'd51547: out <= 16'h0327;
    16'd51548: out <= 16'h0197;    16'd51549: out <= 16'h00FF;    16'd51550: out <= 16'h0211;    16'd51551: out <= 16'h06C4;
    16'd51552: out <= 16'h04E2;    16'd51553: out <= 16'h03FC;    16'd51554: out <= 16'h0435;    16'd51555: out <= 16'hFF0C;
    16'd51556: out <= 16'h0932;    16'd51557: out <= 16'h0130;    16'd51558: out <= 16'h04E0;    16'd51559: out <= 16'h0593;
    16'd51560: out <= 16'h0166;    16'd51561: out <= 16'h00CD;    16'd51562: out <= 16'hFC3C;    16'd51563: out <= 16'hFCDB;
    16'd51564: out <= 16'h0234;    16'd51565: out <= 16'hFBDF;    16'd51566: out <= 16'h017A;    16'd51567: out <= 16'hF758;
    16'd51568: out <= 16'hFD00;    16'd51569: out <= 16'h0676;    16'd51570: out <= 16'h0324;    16'd51571: out <= 16'hFB72;
    16'd51572: out <= 16'h0783;    16'd51573: out <= 16'hFC02;    16'd51574: out <= 16'h04B2;    16'd51575: out <= 16'hFE5D;
    16'd51576: out <= 16'hFB2A;    16'd51577: out <= 16'h01DC;    16'd51578: out <= 16'h0106;    16'd51579: out <= 16'h02A5;
    16'd51580: out <= 16'h00C3;    16'd51581: out <= 16'h002B;    16'd51582: out <= 16'h04DB;    16'd51583: out <= 16'h0AAF;
    16'd51584: out <= 16'h0221;    16'd51585: out <= 16'h0BCF;    16'd51586: out <= 16'h0749;    16'd51587: out <= 16'h0060;
    16'd51588: out <= 16'h045E;    16'd51589: out <= 16'h067F;    16'd51590: out <= 16'h0162;    16'd51591: out <= 16'h01DD;
    16'd51592: out <= 16'h02DD;    16'd51593: out <= 16'hFF4F;    16'd51594: out <= 16'h03CA;    16'd51595: out <= 16'hFF61;
    16'd51596: out <= 16'h049F;    16'd51597: out <= 16'h0079;    16'd51598: out <= 16'h08CC;    16'd51599: out <= 16'hF9FD;
    16'd51600: out <= 16'h0487;    16'd51601: out <= 16'h01BE;    16'd51602: out <= 16'h023C;    16'd51603: out <= 16'h06AE;
    16'd51604: out <= 16'h058E;    16'd51605: out <= 16'h069E;    16'd51606: out <= 16'hFEC0;    16'd51607: out <= 16'h0089;
    16'd51608: out <= 16'h03FF;    16'd51609: out <= 16'h041F;    16'd51610: out <= 16'h061A;    16'd51611: out <= 16'h0400;
    16'd51612: out <= 16'h06D6;    16'd51613: out <= 16'hFDF6;    16'd51614: out <= 16'h0104;    16'd51615: out <= 16'h01B2;
    16'd51616: out <= 16'hFFF1;    16'd51617: out <= 16'h0426;    16'd51618: out <= 16'h0B15;    16'd51619: out <= 16'h0352;
    16'd51620: out <= 16'hFF13;    16'd51621: out <= 16'h046A;    16'd51622: out <= 16'hFF79;    16'd51623: out <= 16'h0455;
    16'd51624: out <= 16'h0222;    16'd51625: out <= 16'h000B;    16'd51626: out <= 16'h0475;    16'd51627: out <= 16'h03CA;
    16'd51628: out <= 16'h0757;    16'd51629: out <= 16'h04AB;    16'd51630: out <= 16'h0733;    16'd51631: out <= 16'h00CA;
    16'd51632: out <= 16'h0BBF;    16'd51633: out <= 16'h0B01;    16'd51634: out <= 16'hFFAC;    16'd51635: out <= 16'h0384;
    16'd51636: out <= 16'hFF1F;    16'd51637: out <= 16'h0361;    16'd51638: out <= 16'h05B4;    16'd51639: out <= 16'h0987;
    16'd51640: out <= 16'h0A55;    16'd51641: out <= 16'h0099;    16'd51642: out <= 16'h00F3;    16'd51643: out <= 16'h013B;
    16'd51644: out <= 16'h0556;    16'd51645: out <= 16'h03DF;    16'd51646: out <= 16'h02FE;    16'd51647: out <= 16'hFEFC;
    16'd51648: out <= 16'hFD88;    16'd51649: out <= 16'hFE0A;    16'd51650: out <= 16'hFE13;    16'd51651: out <= 16'h0043;
    16'd51652: out <= 16'h0246;    16'd51653: out <= 16'hFED4;    16'd51654: out <= 16'h05A6;    16'd51655: out <= 16'hFCFE;
    16'd51656: out <= 16'h095D;    16'd51657: out <= 16'hFC3B;    16'd51658: out <= 16'hFF76;    16'd51659: out <= 16'hFE7C;
    16'd51660: out <= 16'h0531;    16'd51661: out <= 16'hF933;    16'd51662: out <= 16'h0188;    16'd51663: out <= 16'hFDE5;
    16'd51664: out <= 16'h02E0;    16'd51665: out <= 16'h0383;    16'd51666: out <= 16'h0810;    16'd51667: out <= 16'h0A7A;
    16'd51668: out <= 16'hFF06;    16'd51669: out <= 16'hFF21;    16'd51670: out <= 16'hFFEB;    16'd51671: out <= 16'hFFAF;
    16'd51672: out <= 16'h016D;    16'd51673: out <= 16'hFCF3;    16'd51674: out <= 16'hFD8C;    16'd51675: out <= 16'h032B;
    16'd51676: out <= 16'h05AC;    16'd51677: out <= 16'hFE54;    16'd51678: out <= 16'hFB93;    16'd51679: out <= 16'h0543;
    16'd51680: out <= 16'hFDD3;    16'd51681: out <= 16'h021A;    16'd51682: out <= 16'hFD44;    16'd51683: out <= 16'hF95C;
    16'd51684: out <= 16'h02BE;    16'd51685: out <= 16'hFB0C;    16'd51686: out <= 16'h04B7;    16'd51687: out <= 16'h0304;
    16'd51688: out <= 16'hFFC0;    16'd51689: out <= 16'h00A6;    16'd51690: out <= 16'hF9E3;    16'd51691: out <= 16'h0309;
    16'd51692: out <= 16'hFA59;    16'd51693: out <= 16'hFEA9;    16'd51694: out <= 16'h03DF;    16'd51695: out <= 16'hF9F8;
    16'd51696: out <= 16'hF70D;    16'd51697: out <= 16'h0084;    16'd51698: out <= 16'h06A1;    16'd51699: out <= 16'h0037;
    16'd51700: out <= 16'h0049;    16'd51701: out <= 16'hF440;    16'd51702: out <= 16'hFE7E;    16'd51703: out <= 16'h0314;
    16'd51704: out <= 16'hFF6B;    16'd51705: out <= 16'h013F;    16'd51706: out <= 16'hFD04;    16'd51707: out <= 16'h0648;
    16'd51708: out <= 16'hFEB1;    16'd51709: out <= 16'hFB00;    16'd51710: out <= 16'hFD3F;    16'd51711: out <= 16'h007F;
    16'd51712: out <= 16'h0469;    16'd51713: out <= 16'h01A7;    16'd51714: out <= 16'h0672;    16'd51715: out <= 16'h07F4;
    16'd51716: out <= 16'h0113;    16'd51717: out <= 16'h0507;    16'd51718: out <= 16'hFA1C;    16'd51719: out <= 16'h00BD;
    16'd51720: out <= 16'hFF16;    16'd51721: out <= 16'hF6C2;    16'd51722: out <= 16'hFE3A;    16'd51723: out <= 16'h01A0;
    16'd51724: out <= 16'h020A;    16'd51725: out <= 16'h00CA;    16'd51726: out <= 16'h083F;    16'd51727: out <= 16'hF9E2;
    16'd51728: out <= 16'hFB9A;    16'd51729: out <= 16'hFC08;    16'd51730: out <= 16'h0037;    16'd51731: out <= 16'h04BA;
    16'd51732: out <= 16'hF8C6;    16'd51733: out <= 16'h02EE;    16'd51734: out <= 16'hF8E8;    16'd51735: out <= 16'hFE6D;
    16'd51736: out <= 16'hF9B3;    16'd51737: out <= 16'h01A3;    16'd51738: out <= 16'h0177;    16'd51739: out <= 16'h0188;
    16'd51740: out <= 16'hF6AB;    16'd51741: out <= 16'hF9EC;    16'd51742: out <= 16'hFE6F;    16'd51743: out <= 16'hF7FA;
    16'd51744: out <= 16'hF864;    16'd51745: out <= 16'h001D;    16'd51746: out <= 16'h03BF;    16'd51747: out <= 16'h02C9;
    16'd51748: out <= 16'hFBA2;    16'd51749: out <= 16'h052A;    16'd51750: out <= 16'hFD7E;    16'd51751: out <= 16'h06CE;
    16'd51752: out <= 16'h01D3;    16'd51753: out <= 16'hFDE1;    16'd51754: out <= 16'hFF7E;    16'd51755: out <= 16'h01A7;
    16'd51756: out <= 16'hFBE2;    16'd51757: out <= 16'h085B;    16'd51758: out <= 16'h0017;    16'd51759: out <= 16'h0104;
    16'd51760: out <= 16'h0973;    16'd51761: out <= 16'hFE27;    16'd51762: out <= 16'h016C;    16'd51763: out <= 16'h02AD;
    16'd51764: out <= 16'h0250;    16'd51765: out <= 16'h030C;    16'd51766: out <= 16'hFCED;    16'd51767: out <= 16'h0146;
    16'd51768: out <= 16'h01BF;    16'd51769: out <= 16'h03C8;    16'd51770: out <= 16'h0017;    16'd51771: out <= 16'h0368;
    16'd51772: out <= 16'h085C;    16'd51773: out <= 16'h0197;    16'd51774: out <= 16'h0131;    16'd51775: out <= 16'h02CB;
    16'd51776: out <= 16'h00DD;    16'd51777: out <= 16'hFC9D;    16'd51778: out <= 16'hFF06;    16'd51779: out <= 16'h04E9;
    16'd51780: out <= 16'h0173;    16'd51781: out <= 16'hFDCA;    16'd51782: out <= 16'h079A;    16'd51783: out <= 16'hFFAD;
    16'd51784: out <= 16'h0221;    16'd51785: out <= 16'h0452;    16'd51786: out <= 16'h01E3;    16'd51787: out <= 16'h0531;
    16'd51788: out <= 16'h0347;    16'd51789: out <= 16'h0623;    16'd51790: out <= 16'h0491;    16'd51791: out <= 16'h07C7;
    16'd51792: out <= 16'h04B3;    16'd51793: out <= 16'h03C0;    16'd51794: out <= 16'h07DA;    16'd51795: out <= 16'h0773;
    16'd51796: out <= 16'h0437;    16'd51797: out <= 16'h021B;    16'd51798: out <= 16'h043E;    16'd51799: out <= 16'h053C;
    16'd51800: out <= 16'h011B;    16'd51801: out <= 16'h087D;    16'd51802: out <= 16'h0853;    16'd51803: out <= 16'h03AB;
    16'd51804: out <= 16'h0978;    16'd51805: out <= 16'h07D8;    16'd51806: out <= 16'h024A;    16'd51807: out <= 16'h072A;
    16'd51808: out <= 16'h0CAC;    16'd51809: out <= 16'hFEC8;    16'd51810: out <= 16'h0273;    16'd51811: out <= 16'hFFDB;
    16'd51812: out <= 16'h0715;    16'd51813: out <= 16'h0387;    16'd51814: out <= 16'h080D;    16'd51815: out <= 16'hFC0E;
    16'd51816: out <= 16'h04E8;    16'd51817: out <= 16'hFF03;    16'd51818: out <= 16'hFB8E;    16'd51819: out <= 16'h03F0;
    16'd51820: out <= 16'h03B3;    16'd51821: out <= 16'hFCC9;    16'd51822: out <= 16'h01E7;    16'd51823: out <= 16'h0558;
    16'd51824: out <= 16'h048E;    16'd51825: out <= 16'h0138;    16'd51826: out <= 16'h047A;    16'd51827: out <= 16'h027B;
    16'd51828: out <= 16'hFE0F;    16'd51829: out <= 16'h0217;    16'd51830: out <= 16'h06C8;    16'd51831: out <= 16'h01A6;
    16'd51832: out <= 16'h0279;    16'd51833: out <= 16'hFFC7;    16'd51834: out <= 16'hFF78;    16'd51835: out <= 16'h0290;
    16'd51836: out <= 16'h0072;    16'd51837: out <= 16'hFFD9;    16'd51838: out <= 16'h036F;    16'd51839: out <= 16'h06C5;
    16'd51840: out <= 16'h0A7A;    16'd51841: out <= 16'h0BFB;    16'd51842: out <= 16'h007B;    16'd51843: out <= 16'h078E;
    16'd51844: out <= 16'h01DA;    16'd51845: out <= 16'h0535;    16'd51846: out <= 16'h048E;    16'd51847: out <= 16'h069B;
    16'd51848: out <= 16'h026F;    16'd51849: out <= 16'h0525;    16'd51850: out <= 16'hFBB5;    16'd51851: out <= 16'h0124;
    16'd51852: out <= 16'h0260;    16'd51853: out <= 16'h04CC;    16'd51854: out <= 16'h08EA;    16'd51855: out <= 16'h031A;
    16'd51856: out <= 16'h0584;    16'd51857: out <= 16'h0962;    16'd51858: out <= 16'h0925;    16'd51859: out <= 16'h0115;
    16'd51860: out <= 16'h0617;    16'd51861: out <= 16'h000E;    16'd51862: out <= 16'h0643;    16'd51863: out <= 16'h0414;
    16'd51864: out <= 16'hFF4C;    16'd51865: out <= 16'hFF9D;    16'd51866: out <= 16'h0504;    16'd51867: out <= 16'h050D;
    16'd51868: out <= 16'h0681;    16'd51869: out <= 16'hFED2;    16'd51870: out <= 16'h04C0;    16'd51871: out <= 16'h05AA;
    16'd51872: out <= 16'h0609;    16'd51873: out <= 16'h041F;    16'd51874: out <= 16'hFD30;    16'd51875: out <= 16'hFFB8;
    16'd51876: out <= 16'h05BF;    16'd51877: out <= 16'h0257;    16'd51878: out <= 16'hFE4E;    16'd51879: out <= 16'h024D;
    16'd51880: out <= 16'h057C;    16'd51881: out <= 16'h0810;    16'd51882: out <= 16'h0577;    16'd51883: out <= 16'h0B89;
    16'd51884: out <= 16'h0749;    16'd51885: out <= 16'hFFF7;    16'd51886: out <= 16'h0520;    16'd51887: out <= 16'h0932;
    16'd51888: out <= 16'h03DE;    16'd51889: out <= 16'hFC1D;    16'd51890: out <= 16'h0695;    16'd51891: out <= 16'h09AC;
    16'd51892: out <= 16'h0107;    16'd51893: out <= 16'h0304;    16'd51894: out <= 16'h0208;    16'd51895: out <= 16'h066B;
    16'd51896: out <= 16'h0BCE;    16'd51897: out <= 16'h02E5;    16'd51898: out <= 16'h009C;    16'd51899: out <= 16'h02F4;
    16'd51900: out <= 16'h0A5A;    16'd51901: out <= 16'h020A;    16'd51902: out <= 16'hFC5E;    16'd51903: out <= 16'h078E;
    16'd51904: out <= 16'h07B7;    16'd51905: out <= 16'h0870;    16'd51906: out <= 16'h05F0;    16'd51907: out <= 16'h0036;
    16'd51908: out <= 16'hF9BA;    16'd51909: out <= 16'hFE34;    16'd51910: out <= 16'hFE28;    16'd51911: out <= 16'hFD14;
    16'd51912: out <= 16'hFEAB;    16'd51913: out <= 16'h036A;    16'd51914: out <= 16'h0062;    16'd51915: out <= 16'hFED1;
    16'd51916: out <= 16'hFEF4;    16'd51917: out <= 16'h0326;    16'd51918: out <= 16'h02FC;    16'd51919: out <= 16'h04FA;
    16'd51920: out <= 16'hFF85;    16'd51921: out <= 16'h02E6;    16'd51922: out <= 16'hF8B3;    16'd51923: out <= 16'hFADA;
    16'd51924: out <= 16'hFCBF;    16'd51925: out <= 16'hFAB5;    16'd51926: out <= 16'h0213;    16'd51927: out <= 16'h006D;
    16'd51928: out <= 16'h060F;    16'd51929: out <= 16'hFD9D;    16'd51930: out <= 16'hFB83;    16'd51931: out <= 16'hFDD4;
    16'd51932: out <= 16'hFFD3;    16'd51933: out <= 16'hFF8A;    16'd51934: out <= 16'hFCCD;    16'd51935: out <= 16'hF929;
    16'd51936: out <= 16'hFDAD;    16'd51937: out <= 16'hFAB6;    16'd51938: out <= 16'hFE3D;    16'd51939: out <= 16'h03A3;
    16'd51940: out <= 16'hFC74;    16'd51941: out <= 16'hFE07;    16'd51942: out <= 16'hFA92;    16'd51943: out <= 16'hFE46;
    16'd51944: out <= 16'hFD8E;    16'd51945: out <= 16'h022C;    16'd51946: out <= 16'h00EA;    16'd51947: out <= 16'hFA30;
    16'd51948: out <= 16'h05E9;    16'd51949: out <= 16'h0350;    16'd51950: out <= 16'h041D;    16'd51951: out <= 16'h002E;
    16'd51952: out <= 16'hFCEA;    16'd51953: out <= 16'hF67F;    16'd51954: out <= 16'h0169;    16'd51955: out <= 16'hFBBB;
    16'd51956: out <= 16'h007F;    16'd51957: out <= 16'hFBEA;    16'd51958: out <= 16'hFEE9;    16'd51959: out <= 16'hFC03;
    16'd51960: out <= 16'hFEF0;    16'd51961: out <= 16'h02C3;    16'd51962: out <= 16'h05F5;    16'd51963: out <= 16'h0097;
    16'd51964: out <= 16'hFFC6;    16'd51965: out <= 16'h065F;    16'd51966: out <= 16'h0765;    16'd51967: out <= 16'h01A6;
    16'd51968: out <= 16'hFEBB;    16'd51969: out <= 16'h02D5;    16'd51970: out <= 16'hFDCA;    16'd51971: out <= 16'hFE28;
    16'd51972: out <= 16'h00AF;    16'd51973: out <= 16'h0444;    16'd51974: out <= 16'h005B;    16'd51975: out <= 16'h06A9;
    16'd51976: out <= 16'hFB19;    16'd51977: out <= 16'h0375;    16'd51978: out <= 16'hFD80;    16'd51979: out <= 16'hFBB8;
    16'd51980: out <= 16'h02ED;    16'd51981: out <= 16'hFC28;    16'd51982: out <= 16'h017F;    16'd51983: out <= 16'h04BC;
    16'd51984: out <= 16'h04B9;    16'd51985: out <= 16'hFC8A;    16'd51986: out <= 16'hFE24;    16'd51987: out <= 16'hFFFE;
    16'd51988: out <= 16'hFBF1;    16'd51989: out <= 16'h02D1;    16'd51990: out <= 16'hFFA7;    16'd51991: out <= 16'h0147;
    16'd51992: out <= 16'hFBDD;    16'd51993: out <= 16'hF9EC;    16'd51994: out <= 16'hFC39;    16'd51995: out <= 16'h01E7;
    16'd51996: out <= 16'h0559;    16'd51997: out <= 16'h03D6;    16'd51998: out <= 16'h0077;    16'd51999: out <= 16'h0305;
    16'd52000: out <= 16'h00BB;    16'd52001: out <= 16'h01D3;    16'd52002: out <= 16'h0339;    16'd52003: out <= 16'hFD70;
    16'd52004: out <= 16'h062C;    16'd52005: out <= 16'hFB87;    16'd52006: out <= 16'h002D;    16'd52007: out <= 16'h006E;
    16'd52008: out <= 16'hFBFD;    16'd52009: out <= 16'hFC43;    16'd52010: out <= 16'hF72A;    16'd52011: out <= 16'hFDF4;
    16'd52012: out <= 16'h02C5;    16'd52013: out <= 16'h0435;    16'd52014: out <= 16'h0AC2;    16'd52015: out <= 16'hFE61;
    16'd52016: out <= 16'h0140;    16'd52017: out <= 16'h0A94;    16'd52018: out <= 16'h025D;    16'd52019: out <= 16'h0B26;
    16'd52020: out <= 16'h022C;    16'd52021: out <= 16'h0521;    16'd52022: out <= 16'h03CA;    16'd52023: out <= 16'h063C;
    16'd52024: out <= 16'h0261;    16'd52025: out <= 16'h06EC;    16'd52026: out <= 16'h0535;    16'd52027: out <= 16'h06D2;
    16'd52028: out <= 16'hF95C;    16'd52029: out <= 16'h048B;    16'd52030: out <= 16'h04F4;    16'd52031: out <= 16'h0637;
    16'd52032: out <= 16'h0641;    16'd52033: out <= 16'h01A8;    16'd52034: out <= 16'hFBA5;    16'd52035: out <= 16'h01E7;
    16'd52036: out <= 16'h0A14;    16'd52037: out <= 16'h02A0;    16'd52038: out <= 16'h02A9;    16'd52039: out <= 16'h0443;
    16'd52040: out <= 16'h0411;    16'd52041: out <= 16'h071A;    16'd52042: out <= 16'h022D;    16'd52043: out <= 16'h0434;
    16'd52044: out <= 16'h02F6;    16'd52045: out <= 16'h083A;    16'd52046: out <= 16'h0043;    16'd52047: out <= 16'h0B2C;
    16'd52048: out <= 16'h05C5;    16'd52049: out <= 16'h021B;    16'd52050: out <= 16'h03D6;    16'd52051: out <= 16'hFE09;
    16'd52052: out <= 16'hFFAC;    16'd52053: out <= 16'hFDD0;    16'd52054: out <= 16'h0559;    16'd52055: out <= 16'h0765;
    16'd52056: out <= 16'h07EC;    16'd52057: out <= 16'hFFB4;    16'd52058: out <= 16'h0974;    16'd52059: out <= 16'h049C;
    16'd52060: out <= 16'h071B;    16'd52061: out <= 16'h0426;    16'd52062: out <= 16'h0454;    16'd52063: out <= 16'h08FA;
    16'd52064: out <= 16'h05C1;    16'd52065: out <= 16'h0379;    16'd52066: out <= 16'h00DB;    16'd52067: out <= 16'h04D1;
    16'd52068: out <= 16'hFE1F;    16'd52069: out <= 16'h0485;    16'd52070: out <= 16'h0040;    16'd52071: out <= 16'hF890;
    16'd52072: out <= 16'h0220;    16'd52073: out <= 16'hFE26;    16'd52074: out <= 16'h043B;    16'd52075: out <= 16'hFE01;
    16'd52076: out <= 16'h02C7;    16'd52077: out <= 16'h0298;    16'd52078: out <= 16'h05C7;    16'd52079: out <= 16'hFB83;
    16'd52080: out <= 16'h03A9;    16'd52081: out <= 16'hFF97;    16'd52082: out <= 16'hFD52;    16'd52083: out <= 16'hFAC6;
    16'd52084: out <= 16'hFF42;    16'd52085: out <= 16'hFB88;    16'd52086: out <= 16'h02CA;    16'd52087: out <= 16'hFFAF;
    16'd52088: out <= 16'hFA34;    16'd52089: out <= 16'hFF32;    16'd52090: out <= 16'hFEFC;    16'd52091: out <= 16'hFDA9;
    16'd52092: out <= 16'hFBCE;    16'd52093: out <= 16'hFEFC;    16'd52094: out <= 16'h02C9;    16'd52095: out <= 16'h0B3D;
    16'd52096: out <= 16'h00DC;    16'd52097: out <= 16'h08A9;    16'd52098: out <= 16'h0B46;    16'd52099: out <= 16'h09FB;
    16'd52100: out <= 16'h0311;    16'd52101: out <= 16'h0753;    16'd52102: out <= 16'h0760;    16'd52103: out <= 16'h06E8;
    16'd52104: out <= 16'h0AE2;    16'd52105: out <= 16'h0485;    16'd52106: out <= 16'h02C0;    16'd52107: out <= 16'hFF1A;
    16'd52108: out <= 16'h0415;    16'd52109: out <= 16'hFDFA;    16'd52110: out <= 16'h02F9;    16'd52111: out <= 16'h05A1;
    16'd52112: out <= 16'h0638;    16'd52113: out <= 16'h0706;    16'd52114: out <= 16'h031A;    16'd52115: out <= 16'h01F0;
    16'd52116: out <= 16'hFD4A;    16'd52117: out <= 16'h00B3;    16'd52118: out <= 16'h045D;    16'd52119: out <= 16'h018F;
    16'd52120: out <= 16'h0369;    16'd52121: out <= 16'h06C8;    16'd52122: out <= 16'h02E3;    16'd52123: out <= 16'h0505;
    16'd52124: out <= 16'h00F7;    16'd52125: out <= 16'h02B7;    16'd52126: out <= 16'h0734;    16'd52127: out <= 16'h09A7;
    16'd52128: out <= 16'h0650;    16'd52129: out <= 16'h0576;    16'd52130: out <= 16'h036D;    16'd52131: out <= 16'hFBBA;
    16'd52132: out <= 16'h02F9;    16'd52133: out <= 16'h051A;    16'd52134: out <= 16'h05C5;    16'd52135: out <= 16'h02D6;
    16'd52136: out <= 16'h0088;    16'd52137: out <= 16'hFFE4;    16'd52138: out <= 16'h0705;    16'd52139: out <= 16'h081F;
    16'd52140: out <= 16'h0863;    16'd52141: out <= 16'h00F3;    16'd52142: out <= 16'h09B2;    16'd52143: out <= 16'h051B;
    16'd52144: out <= 16'h043B;    16'd52145: out <= 16'h08ED;    16'd52146: out <= 16'h0561;    16'd52147: out <= 16'h0439;
    16'd52148: out <= 16'h05DA;    16'd52149: out <= 16'h0481;    16'd52150: out <= 16'h0460;    16'd52151: out <= 16'h036D;
    16'd52152: out <= 16'h03EF;    16'd52153: out <= 16'hFFCF;    16'd52154: out <= 16'hFE4A;    16'd52155: out <= 16'h0342;
    16'd52156: out <= 16'h02EA;    16'd52157: out <= 16'h0621;    16'd52158: out <= 16'h06F7;    16'd52159: out <= 16'h057E;
    16'd52160: out <= 16'h029D;    16'd52161: out <= 16'h0414;    16'd52162: out <= 16'h014A;    16'd52163: out <= 16'h0530;
    16'd52164: out <= 16'hFB6D;    16'd52165: out <= 16'hFF53;    16'd52166: out <= 16'hFFED;    16'd52167: out <= 16'h049B;
    16'd52168: out <= 16'h0503;    16'd52169: out <= 16'h0328;    16'd52170: out <= 16'h052A;    16'd52171: out <= 16'hF712;
    16'd52172: out <= 16'h025C;    16'd52173: out <= 16'hFE27;    16'd52174: out <= 16'h00F7;    16'd52175: out <= 16'h0264;
    16'd52176: out <= 16'hFACA;    16'd52177: out <= 16'h007E;    16'd52178: out <= 16'h01E3;    16'd52179: out <= 16'h02F3;
    16'd52180: out <= 16'h0358;    16'd52181: out <= 16'hF572;    16'd52182: out <= 16'hFE47;    16'd52183: out <= 16'h008C;
    16'd52184: out <= 16'h06A3;    16'd52185: out <= 16'hF92A;    16'd52186: out <= 16'hFC86;    16'd52187: out <= 16'hF63C;
    16'd52188: out <= 16'h03D5;    16'd52189: out <= 16'hFC9B;    16'd52190: out <= 16'h02EE;    16'd52191: out <= 16'h00E0;
    16'd52192: out <= 16'hFF54;    16'd52193: out <= 16'h01B4;    16'd52194: out <= 16'hFC2C;    16'd52195: out <= 16'h0486;
    16'd52196: out <= 16'hF946;    16'd52197: out <= 16'hF6F3;    16'd52198: out <= 16'h0041;    16'd52199: out <= 16'h0381;
    16'd52200: out <= 16'hFFAF;    16'd52201: out <= 16'h0168;    16'd52202: out <= 16'h0A97;    16'd52203: out <= 16'hFEBB;
    16'd52204: out <= 16'hFC06;    16'd52205: out <= 16'h01AB;    16'd52206: out <= 16'hFCF4;    16'd52207: out <= 16'h033D;
    16'd52208: out <= 16'h0427;    16'd52209: out <= 16'h00EC;    16'd52210: out <= 16'hFCEC;    16'd52211: out <= 16'h0054;
    16'd52212: out <= 16'h019F;    16'd52213: out <= 16'hFE0A;    16'd52214: out <= 16'hFE8D;    16'd52215: out <= 16'h081F;
    16'd52216: out <= 16'hFC63;    16'd52217: out <= 16'hFD8D;    16'd52218: out <= 16'h011F;    16'd52219: out <= 16'hFD35;
    16'd52220: out <= 16'hFF10;    16'd52221: out <= 16'hFE5D;    16'd52222: out <= 16'h0342;    16'd52223: out <= 16'hFEB3;
    16'd52224: out <= 16'hFCAD;    16'd52225: out <= 16'hFB4D;    16'd52226: out <= 16'h004B;    16'd52227: out <= 16'h005F;
    16'd52228: out <= 16'h02A2;    16'd52229: out <= 16'h02F5;    16'd52230: out <= 16'hFE7B;    16'd52231: out <= 16'hF6D8;
    16'd52232: out <= 16'h0478;    16'd52233: out <= 16'h0409;    16'd52234: out <= 16'hFB57;    16'd52235: out <= 16'h06AF;
    16'd52236: out <= 16'h068A;    16'd52237: out <= 16'h00B4;    16'd52238: out <= 16'h0419;    16'd52239: out <= 16'h0A92;
    16'd52240: out <= 16'h0466;    16'd52241: out <= 16'h01E9;    16'd52242: out <= 16'hFEA9;    16'd52243: out <= 16'hFABE;
    16'd52244: out <= 16'h0543;    16'd52245: out <= 16'h065B;    16'd52246: out <= 16'hFAB7;    16'd52247: out <= 16'hFB79;
    16'd52248: out <= 16'h0699;    16'd52249: out <= 16'h01DF;    16'd52250: out <= 16'hFF7C;    16'd52251: out <= 16'hFCB2;
    16'd52252: out <= 16'h0303;    16'd52253: out <= 16'h0185;    16'd52254: out <= 16'hFC77;    16'd52255: out <= 16'h0162;
    16'd52256: out <= 16'hFD3D;    16'd52257: out <= 16'hFDF8;    16'd52258: out <= 16'hFF34;    16'd52259: out <= 16'h0350;
    16'd52260: out <= 16'hF801;    16'd52261: out <= 16'h02AE;    16'd52262: out <= 16'h04CD;    16'd52263: out <= 16'hFDBD;
    16'd52264: out <= 16'hFC21;    16'd52265: out <= 16'h0694;    16'd52266: out <= 16'hFC67;    16'd52267: out <= 16'h0652;
    16'd52268: out <= 16'h03AA;    16'd52269: out <= 16'h0194;    16'd52270: out <= 16'h002E;    16'd52271: out <= 16'hFE21;
    16'd52272: out <= 16'h06F8;    16'd52273: out <= 16'hFB54;    16'd52274: out <= 16'h04A6;    16'd52275: out <= 16'h06B1;
    16'd52276: out <= 16'h021D;    16'd52277: out <= 16'h0315;    16'd52278: out <= 16'h0E41;    16'd52279: out <= 16'h005B;
    16'd52280: out <= 16'h035D;    16'd52281: out <= 16'h0380;    16'd52282: out <= 16'h0271;    16'd52283: out <= 16'h01C2;
    16'd52284: out <= 16'h0861;    16'd52285: out <= 16'h04A0;    16'd52286: out <= 16'h05A5;    16'd52287: out <= 16'h047D;
    16'd52288: out <= 16'h011F;    16'd52289: out <= 16'h0591;    16'd52290: out <= 16'h0149;    16'd52291: out <= 16'h055D;
    16'd52292: out <= 16'h0AF2;    16'd52293: out <= 16'h0BB6;    16'd52294: out <= 16'h0551;    16'd52295: out <= 16'h0A40;
    16'd52296: out <= 16'h0568;    16'd52297: out <= 16'hFAE4;    16'd52298: out <= 16'h04C6;    16'd52299: out <= 16'h06B2;
    16'd52300: out <= 16'h0651;    16'd52301: out <= 16'h04CF;    16'd52302: out <= 16'h0837;    16'd52303: out <= 16'h0347;
    16'd52304: out <= 16'h00A6;    16'd52305: out <= 16'h0717;    16'd52306: out <= 16'h007F;    16'd52307: out <= 16'h06CA;
    16'd52308: out <= 16'h05AB;    16'd52309: out <= 16'h00F8;    16'd52310: out <= 16'h001B;    16'd52311: out <= 16'h0801;
    16'd52312: out <= 16'h02C3;    16'd52313: out <= 16'h0089;    16'd52314: out <= 16'h0751;    16'd52315: out <= 16'h0473;
    16'd52316: out <= 16'h0237;    16'd52317: out <= 16'h028C;    16'd52318: out <= 16'h05CB;    16'd52319: out <= 16'h083C;
    16'd52320: out <= 16'h0791;    16'd52321: out <= 16'h0091;    16'd52322: out <= 16'h0018;    16'd52323: out <= 16'hFF65;
    16'd52324: out <= 16'h04E1;    16'd52325: out <= 16'hFD2D;    16'd52326: out <= 16'hFBBF;    16'd52327: out <= 16'h0A38;
    16'd52328: out <= 16'h015C;    16'd52329: out <= 16'h0360;    16'd52330: out <= 16'hFB14;    16'd52331: out <= 16'hFE7F;
    16'd52332: out <= 16'hFB8C;    16'd52333: out <= 16'hFEDF;    16'd52334: out <= 16'hFE2E;    16'd52335: out <= 16'h03FC;
    16'd52336: out <= 16'hFC74;    16'd52337: out <= 16'hFBAF;    16'd52338: out <= 16'hFA24;    16'd52339: out <= 16'h0370;
    16'd52340: out <= 16'h0002;    16'd52341: out <= 16'hFC99;    16'd52342: out <= 16'h0220;    16'd52343: out <= 16'hFE83;
    16'd52344: out <= 16'h01A1;    16'd52345: out <= 16'h034F;    16'd52346: out <= 16'hFDBA;    16'd52347: out <= 16'hFC8F;
    16'd52348: out <= 16'h057D;    16'd52349: out <= 16'h02CC;    16'd52350: out <= 16'hFAEA;    16'd52351: out <= 16'hFFC3;
    16'd52352: out <= 16'h026A;    16'd52353: out <= 16'h05A6;    16'd52354: out <= 16'h05C2;    16'd52355: out <= 16'h03FF;
    16'd52356: out <= 16'h0646;    16'd52357: out <= 16'h04B5;    16'd52358: out <= 16'hFD2A;    16'd52359: out <= 16'h031A;
    16'd52360: out <= 16'h049D;    16'd52361: out <= 16'hF89E;    16'd52362: out <= 16'h01E5;    16'd52363: out <= 16'h0277;
    16'd52364: out <= 16'hFF2F;    16'd52365: out <= 16'h08F9;    16'd52366: out <= 16'h05C8;    16'd52367: out <= 16'h0525;
    16'd52368: out <= 16'h0918;    16'd52369: out <= 16'h02FF;    16'd52370: out <= 16'h07AF;    16'd52371: out <= 16'h0BF5;
    16'd52372: out <= 16'h03B0;    16'd52373: out <= 16'h05E8;    16'd52374: out <= 16'h08D5;    16'd52375: out <= 16'hFEE3;
    16'd52376: out <= 16'h01E0;    16'd52377: out <= 16'hFDD3;    16'd52378: out <= 16'h01CF;    16'd52379: out <= 16'h096B;
    16'd52380: out <= 16'hFDD3;    16'd52381: out <= 16'h066B;    16'd52382: out <= 16'h07A5;    16'd52383: out <= 16'h0517;
    16'd52384: out <= 16'hFD7F;    16'd52385: out <= 16'h04E2;    16'd52386: out <= 16'h0435;    16'd52387: out <= 16'h013F;
    16'd52388: out <= 16'h059D;    16'd52389: out <= 16'h05FB;    16'd52390: out <= 16'h0B8A;    16'd52391: out <= 16'hFFCD;
    16'd52392: out <= 16'h028E;    16'd52393: out <= 16'h01F3;    16'd52394: out <= 16'h03A2;    16'd52395: out <= 16'h054D;
    16'd52396: out <= 16'h03C7;    16'd52397: out <= 16'h08B8;    16'd52398: out <= 16'h03D7;    16'd52399: out <= 16'h0892;
    16'd52400: out <= 16'h0818;    16'd52401: out <= 16'h04FC;    16'd52402: out <= 16'hFDDC;    16'd52403: out <= 16'h003C;
    16'd52404: out <= 16'h049B;    16'd52405: out <= 16'h0461;    16'd52406: out <= 16'h02A5;    16'd52407: out <= 16'h04FD;
    16'd52408: out <= 16'h0126;    16'd52409: out <= 16'h0533;    16'd52410: out <= 16'h0735;    16'd52411: out <= 16'h01A5;
    16'd52412: out <= 16'h08D5;    16'd52413: out <= 16'h0031;    16'd52414: out <= 16'h06F4;    16'd52415: out <= 16'h0A19;
    16'd52416: out <= 16'h033B;    16'd52417: out <= 16'h031C;    16'd52418: out <= 16'h028E;    16'd52419: out <= 16'hFC18;
    16'd52420: out <= 16'hFD74;    16'd52421: out <= 16'h00B2;    16'd52422: out <= 16'hFC1F;    16'd52423: out <= 16'hFCCB;
    16'd52424: out <= 16'h067D;    16'd52425: out <= 16'h0160;    16'd52426: out <= 16'hFF7B;    16'd52427: out <= 16'h0252;
    16'd52428: out <= 16'h03D5;    16'd52429: out <= 16'h029E;    16'd52430: out <= 16'hFF5E;    16'd52431: out <= 16'h05CA;
    16'd52432: out <= 16'h0531;    16'd52433: out <= 16'hFC94;    16'd52434: out <= 16'hFBA2;    16'd52435: out <= 16'h01CC;
    16'd52436: out <= 16'hFA46;    16'd52437: out <= 16'hFE3E;    16'd52438: out <= 16'hF9F2;    16'd52439: out <= 16'hFE0D;
    16'd52440: out <= 16'h0017;    16'd52441: out <= 16'hFEBF;    16'd52442: out <= 16'h0290;    16'd52443: out <= 16'hFC33;
    16'd52444: out <= 16'hFE52;    16'd52445: out <= 16'h002E;    16'd52446: out <= 16'hFF88;    16'd52447: out <= 16'h0018;
    16'd52448: out <= 16'h0146;    16'd52449: out <= 16'h041D;    16'd52450: out <= 16'h0071;    16'd52451: out <= 16'h05D1;
    16'd52452: out <= 16'hF8C6;    16'd52453: out <= 16'hFF24;    16'd52454: out <= 16'h042C;    16'd52455: out <= 16'h0694;
    16'd52456: out <= 16'h016A;    16'd52457: out <= 16'h0008;    16'd52458: out <= 16'hFE98;    16'd52459: out <= 16'hFBFF;
    16'd52460: out <= 16'h045F;    16'd52461: out <= 16'hFCEE;    16'd52462: out <= 16'hFF43;    16'd52463: out <= 16'hF78C;
    16'd52464: out <= 16'h05B0;    16'd52465: out <= 16'hF979;    16'd52466: out <= 16'hFE5A;    16'd52467: out <= 16'hFAAB;
    16'd52468: out <= 16'hFE7F;    16'd52469: out <= 16'hFF07;    16'd52470: out <= 16'h030D;    16'd52471: out <= 16'hF924;
    16'd52472: out <= 16'hFE1B;    16'd52473: out <= 16'h032F;    16'd52474: out <= 16'hFDC9;    16'd52475: out <= 16'h0174;
    16'd52476: out <= 16'h0042;    16'd52477: out <= 16'hF980;    16'd52478: out <= 16'hFCF8;    16'd52479: out <= 16'h01EB;
    16'd52480: out <= 16'h0178;    16'd52481: out <= 16'hFA02;    16'd52482: out <= 16'hFF80;    16'd52483: out <= 16'hFC79;
    16'd52484: out <= 16'hFCA6;    16'd52485: out <= 16'h02DD;    16'd52486: out <= 16'hFE08;    16'd52487: out <= 16'hFC02;
    16'd52488: out <= 16'hFEF5;    16'd52489: out <= 16'h0534;    16'd52490: out <= 16'hF9F2;    16'd52491: out <= 16'h0187;
    16'd52492: out <= 16'h04E1;    16'd52493: out <= 16'h02E8;    16'd52494: out <= 16'h028B;    16'd52495: out <= 16'hFD7D;
    16'd52496: out <= 16'hFF16;    16'd52497: out <= 16'h0047;    16'd52498: out <= 16'h0096;    16'd52499: out <= 16'hF94E;
    16'd52500: out <= 16'hFBA8;    16'd52501: out <= 16'h015A;    16'd52502: out <= 16'hFDDF;    16'd52503: out <= 16'hFD88;
    16'd52504: out <= 16'hFEBF;    16'd52505: out <= 16'h0168;    16'd52506: out <= 16'h002F;    16'd52507: out <= 16'h0225;
    16'd52508: out <= 16'hFBB5;    16'd52509: out <= 16'hFDFC;    16'd52510: out <= 16'hFF07;    16'd52511: out <= 16'hFC32;
    16'd52512: out <= 16'h012D;    16'd52513: out <= 16'h0C7B;    16'd52514: out <= 16'h02E2;    16'd52515: out <= 16'hFFEE;
    16'd52516: out <= 16'h024C;    16'd52517: out <= 16'h03CF;    16'd52518: out <= 16'hF947;    16'd52519: out <= 16'h0388;
    16'd52520: out <= 16'hFD99;    16'd52521: out <= 16'hFBD5;    16'd52522: out <= 16'hFA22;    16'd52523: out <= 16'hFEB5;
    16'd52524: out <= 16'hFBA1;    16'd52525: out <= 16'hFD88;    16'd52526: out <= 16'hFD69;    16'd52527: out <= 16'h0005;
    16'd52528: out <= 16'h0324;    16'd52529: out <= 16'h04E1;    16'd52530: out <= 16'h0661;    16'd52531: out <= 16'h0145;
    16'd52532: out <= 16'h04A1;    16'd52533: out <= 16'h092F;    16'd52534: out <= 16'h0099;    16'd52535: out <= 16'h070C;
    16'd52536: out <= 16'h03D7;    16'd52537: out <= 16'h0557;    16'd52538: out <= 16'h07A7;    16'd52539: out <= 16'h02E2;
    16'd52540: out <= 16'h0BAC;    16'd52541: out <= 16'h0389;    16'd52542: out <= 16'h07FF;    16'd52543: out <= 16'h011B;
    16'd52544: out <= 16'h0332;    16'd52545: out <= 16'h0E8C;    16'd52546: out <= 16'h0848;    16'd52547: out <= 16'h0113;
    16'd52548: out <= 16'h04A1;    16'd52549: out <= 16'h04D9;    16'd52550: out <= 16'h00FB;    16'd52551: out <= 16'h035F;
    16'd52552: out <= 16'hFE94;    16'd52553: out <= 16'h05A7;    16'd52554: out <= 16'h07C5;    16'd52555: out <= 16'h0108;
    16'd52556: out <= 16'h01AD;    16'd52557: out <= 16'hFF74;    16'd52558: out <= 16'h0174;    16'd52559: out <= 16'h0868;
    16'd52560: out <= 16'h079F;    16'd52561: out <= 16'hFECE;    16'd52562: out <= 16'h06DA;    16'd52563: out <= 16'h0179;
    16'd52564: out <= 16'h07A3;    16'd52565: out <= 16'h08AB;    16'd52566: out <= 16'h076E;    16'd52567: out <= 16'h0330;
    16'd52568: out <= 16'h0156;    16'd52569: out <= 16'h013C;    16'd52570: out <= 16'h054E;    16'd52571: out <= 16'h0376;
    16'd52572: out <= 16'h061E;    16'd52573: out <= 16'h06F6;    16'd52574: out <= 16'h0285;    16'd52575: out <= 16'h0AE0;
    16'd52576: out <= 16'h052C;    16'd52577: out <= 16'h0050;    16'd52578: out <= 16'h0375;    16'd52579: out <= 16'hFD4E;
    16'd52580: out <= 16'hFA67;    16'd52581: out <= 16'hFEAF;    16'd52582: out <= 16'h004D;    16'd52583: out <= 16'hF9AE;
    16'd52584: out <= 16'hFC5C;    16'd52585: out <= 16'hFD76;    16'd52586: out <= 16'h05E1;    16'd52587: out <= 16'h07C1;
    16'd52588: out <= 16'hFE3F;    16'd52589: out <= 16'hFDE9;    16'd52590: out <= 16'h0086;    16'd52591: out <= 16'h0441;
    16'd52592: out <= 16'hFCAA;    16'd52593: out <= 16'h011A;    16'd52594: out <= 16'hFABE;    16'd52595: out <= 16'h01F5;
    16'd52596: out <= 16'h05D9;    16'd52597: out <= 16'hFCBE;    16'd52598: out <= 16'h049A;    16'd52599: out <= 16'h002A;
    16'd52600: out <= 16'hFBFD;    16'd52601: out <= 16'hFCBB;    16'd52602: out <= 16'hFF89;    16'd52603: out <= 16'hFC9D;
    16'd52604: out <= 16'h0568;    16'd52605: out <= 16'hFD3E;    16'd52606: out <= 16'h02DF;    16'd52607: out <= 16'hF6EC;
    16'd52608: out <= 16'h0612;    16'd52609: out <= 16'h03DA;    16'd52610: out <= 16'h090D;    16'd52611: out <= 16'hFEEF;
    16'd52612: out <= 16'h003F;    16'd52613: out <= 16'h0FFE;    16'd52614: out <= 16'h034B;    16'd52615: out <= 16'h0549;
    16'd52616: out <= 16'h04EC;    16'd52617: out <= 16'h03CF;    16'd52618: out <= 16'h014B;    16'd52619: out <= 16'hFF24;
    16'd52620: out <= 16'h03E5;    16'd52621: out <= 16'h04F1;    16'd52622: out <= 16'h01FC;    16'd52623: out <= 16'h0BF9;
    16'd52624: out <= 16'h0358;    16'd52625: out <= 16'h05D9;    16'd52626: out <= 16'h0415;    16'd52627: out <= 16'h01F5;
    16'd52628: out <= 16'h034D;    16'd52629: out <= 16'h007C;    16'd52630: out <= 16'h0290;    16'd52631: out <= 16'h000F;
    16'd52632: out <= 16'h01A5;    16'd52633: out <= 16'h0593;    16'd52634: out <= 16'h033B;    16'd52635: out <= 16'h021C;
    16'd52636: out <= 16'h081E;    16'd52637: out <= 16'h035A;    16'd52638: out <= 16'h0450;    16'd52639: out <= 16'h0AC8;
    16'd52640: out <= 16'h0547;    16'd52641: out <= 16'h0602;    16'd52642: out <= 16'hFF38;    16'd52643: out <= 16'h00BC;
    16'd52644: out <= 16'h07AA;    16'd52645: out <= 16'h02CE;    16'd52646: out <= 16'h023C;    16'd52647: out <= 16'h0497;
    16'd52648: out <= 16'h07A1;    16'd52649: out <= 16'h0439;    16'd52650: out <= 16'h08AE;    16'd52651: out <= 16'h0B34;
    16'd52652: out <= 16'h03C3;    16'd52653: out <= 16'h03AE;    16'd52654: out <= 16'h03A5;    16'd52655: out <= 16'h005A;
    16'd52656: out <= 16'h03FD;    16'd52657: out <= 16'h08DE;    16'd52658: out <= 16'h0809;    16'd52659: out <= 16'h0979;
    16'd52660: out <= 16'h041B;    16'd52661: out <= 16'h0A51;    16'd52662: out <= 16'h00EA;    16'd52663: out <= 16'h03C9;
    16'd52664: out <= 16'h0471;    16'd52665: out <= 16'h00BD;    16'd52666: out <= 16'hFEE3;    16'd52667: out <= 16'h06BB;
    16'd52668: out <= 16'h0C15;    16'd52669: out <= 16'hFF07;    16'd52670: out <= 16'h0BBD;    16'd52671: out <= 16'h0756;
    16'd52672: out <= 16'h075D;    16'd52673: out <= 16'h0A48;    16'd52674: out <= 16'h09BD;    16'd52675: out <= 16'hFF38;
    16'd52676: out <= 16'hFB70;    16'd52677: out <= 16'h0056;    16'd52678: out <= 16'hFCD8;    16'd52679: out <= 16'hFEBB;
    16'd52680: out <= 16'h0210;    16'd52681: out <= 16'hFBEC;    16'd52682: out <= 16'h071C;    16'd52683: out <= 16'h0529;
    16'd52684: out <= 16'hFE54;    16'd52685: out <= 16'hFA75;    16'd52686: out <= 16'h011D;    16'd52687: out <= 16'hFA80;
    16'd52688: out <= 16'h01DE;    16'd52689: out <= 16'hFC4A;    16'd52690: out <= 16'h02FE;    16'd52691: out <= 16'hFDDD;
    16'd52692: out <= 16'hFDF9;    16'd52693: out <= 16'hFA02;    16'd52694: out <= 16'h0094;    16'd52695: out <= 16'h019C;
    16'd52696: out <= 16'hFF86;    16'd52697: out <= 16'hFC2E;    16'd52698: out <= 16'h0921;    16'd52699: out <= 16'hFC07;
    16'd52700: out <= 16'hFDB4;    16'd52701: out <= 16'h00BD;    16'd52702: out <= 16'h01C5;    16'd52703: out <= 16'hF7A6;
    16'd52704: out <= 16'h0110;    16'd52705: out <= 16'h00EA;    16'd52706: out <= 16'hFC20;    16'd52707: out <= 16'h04D3;
    16'd52708: out <= 16'h0334;    16'd52709: out <= 16'h03CA;    16'd52710: out <= 16'hFE42;    16'd52711: out <= 16'h0079;
    16'd52712: out <= 16'hFFFD;    16'd52713: out <= 16'h0216;    16'd52714: out <= 16'h05B9;    16'd52715: out <= 16'h061D;
    16'd52716: out <= 16'h0390;    16'd52717: out <= 16'hFAB2;    16'd52718: out <= 16'hF7D6;    16'd52719: out <= 16'hFF4B;
    16'd52720: out <= 16'h0048;    16'd52721: out <= 16'h0103;    16'd52722: out <= 16'h04E4;    16'd52723: out <= 16'hFF81;
    16'd52724: out <= 16'hFF58;    16'd52725: out <= 16'hFFF9;    16'd52726: out <= 16'h020D;    16'd52727: out <= 16'hFCFE;
    16'd52728: out <= 16'hFA62;    16'd52729: out <= 16'h005A;    16'd52730: out <= 16'h0125;    16'd52731: out <= 16'hFDDA;
    16'd52732: out <= 16'hFD71;    16'd52733: out <= 16'h022A;    16'd52734: out <= 16'h02CD;    16'd52735: out <= 16'hFC15;
    16'd52736: out <= 16'h0A8E;    16'd52737: out <= 16'h00C8;    16'd52738: out <= 16'hFFEF;    16'd52739: out <= 16'h02B8;
    16'd52740: out <= 16'h007B;    16'd52741: out <= 16'h02F0;    16'd52742: out <= 16'hFDB4;    16'd52743: out <= 16'hFE09;
    16'd52744: out <= 16'h0127;    16'd52745: out <= 16'hFF91;    16'd52746: out <= 16'hFE13;    16'd52747: out <= 16'hFDEC;
    16'd52748: out <= 16'h00D2;    16'd52749: out <= 16'h01C2;    16'd52750: out <= 16'hFF08;    16'd52751: out <= 16'hFD64;
    16'd52752: out <= 16'h03B2;    16'd52753: out <= 16'h005A;    16'd52754: out <= 16'h02DE;    16'd52755: out <= 16'h016B;
    16'd52756: out <= 16'h025A;    16'd52757: out <= 16'hFC46;    16'd52758: out <= 16'hFFFF;    16'd52759: out <= 16'h0194;
    16'd52760: out <= 16'h0652;    16'd52761: out <= 16'h0448;    16'd52762: out <= 16'h0383;    16'd52763: out <= 16'h0519;
    16'd52764: out <= 16'h0777;    16'd52765: out <= 16'hF79D;    16'd52766: out <= 16'hFB37;    16'd52767: out <= 16'hFE5B;
    16'd52768: out <= 16'h0175;    16'd52769: out <= 16'hFE4F;    16'd52770: out <= 16'h042A;    16'd52771: out <= 16'hFFDE;
    16'd52772: out <= 16'h0761;    16'd52773: out <= 16'hFEBA;    16'd52774: out <= 16'hFD16;    16'd52775: out <= 16'h02D1;
    16'd52776: out <= 16'hFFF8;    16'd52777: out <= 16'hFC39;    16'd52778: out <= 16'hFFF9;    16'd52779: out <= 16'hFEC1;
    16'd52780: out <= 16'hFEA8;    16'd52781: out <= 16'h0292;    16'd52782: out <= 16'h0215;    16'd52783: out <= 16'hF77A;
    16'd52784: out <= 16'h024D;    16'd52785: out <= 16'h0781;    16'd52786: out <= 16'h036C;    16'd52787: out <= 16'h0895;
    16'd52788: out <= 16'h030C;    16'd52789: out <= 16'h05E9;    16'd52790: out <= 16'h062B;    16'd52791: out <= 16'h01C1;
    16'd52792: out <= 16'hFE21;    16'd52793: out <= 16'hFEDB;    16'd52794: out <= 16'h02BD;    16'd52795: out <= 16'h06AF;
    16'd52796: out <= 16'h0873;    16'd52797: out <= 16'h03AA;    16'd52798: out <= 16'h0973;    16'd52799: out <= 16'h012B;
    16'd52800: out <= 16'h04BE;    16'd52801: out <= 16'hFEB5;    16'd52802: out <= 16'h03F2;    16'd52803: out <= 16'h060D;
    16'd52804: out <= 16'h07A3;    16'd52805: out <= 16'hFE38;    16'd52806: out <= 16'h0234;    16'd52807: out <= 16'h0576;
    16'd52808: out <= 16'h02E6;    16'd52809: out <= 16'h022F;    16'd52810: out <= 16'h03DA;    16'd52811: out <= 16'h06B9;
    16'd52812: out <= 16'h07CE;    16'd52813: out <= 16'hFE1B;    16'd52814: out <= 16'h0118;    16'd52815: out <= 16'hFFE3;
    16'd52816: out <= 16'hFCFC;    16'd52817: out <= 16'h0289;    16'd52818: out <= 16'h0709;    16'd52819: out <= 16'h04B1;
    16'd52820: out <= 16'h0454;    16'd52821: out <= 16'h037F;    16'd52822: out <= 16'hFF06;    16'd52823: out <= 16'h049E;
    16'd52824: out <= 16'h0566;    16'd52825: out <= 16'h0122;    16'd52826: out <= 16'hFFBE;    16'd52827: out <= 16'h011B;
    16'd52828: out <= 16'h03B2;    16'd52829: out <= 16'hFF46;    16'd52830: out <= 16'h001E;    16'd52831: out <= 16'h0684;
    16'd52832: out <= 16'hFFD1;    16'd52833: out <= 16'hF7D8;    16'd52834: out <= 16'h0182;    16'd52835: out <= 16'hFC5A;
    16'd52836: out <= 16'hFCF0;    16'd52837: out <= 16'hFE07;    16'd52838: out <= 16'h07AF;    16'd52839: out <= 16'hFF68;
    16'd52840: out <= 16'h059C;    16'd52841: out <= 16'hFC8C;    16'd52842: out <= 16'hFEBF;    16'd52843: out <= 16'h0503;
    16'd52844: out <= 16'h02D0;    16'd52845: out <= 16'hFC2F;    16'd52846: out <= 16'hFE89;    16'd52847: out <= 16'h047B;
    16'd52848: out <= 16'hFC06;    16'd52849: out <= 16'h011C;    16'd52850: out <= 16'hF533;    16'd52851: out <= 16'hFF2D;
    16'd52852: out <= 16'hFC11;    16'd52853: out <= 16'hFA7E;    16'd52854: out <= 16'h02D7;    16'd52855: out <= 16'hFA14;
    16'd52856: out <= 16'h02B1;    16'd52857: out <= 16'hFCFD;    16'd52858: out <= 16'hFD92;    16'd52859: out <= 16'hFF4E;
    16'd52860: out <= 16'hFE55;    16'd52861: out <= 16'h0073;    16'd52862: out <= 16'hFF77;    16'd52863: out <= 16'h0499;
    16'd52864: out <= 16'h06CD;    16'd52865: out <= 16'h0C38;    16'd52866: out <= 16'h000A;    16'd52867: out <= 16'h0713;
    16'd52868: out <= 16'hFFF9;    16'd52869: out <= 16'h0A44;    16'd52870: out <= 16'hFC6E;    16'd52871: out <= 16'h06C7;
    16'd52872: out <= 16'h0906;    16'd52873: out <= 16'h08AC;    16'd52874: out <= 16'h01E5;    16'd52875: out <= 16'h03E1;
    16'd52876: out <= 16'h0121;    16'd52877: out <= 16'h073E;    16'd52878: out <= 16'h03CC;    16'd52879: out <= 16'h09D8;
    16'd52880: out <= 16'h069C;    16'd52881: out <= 16'hFF8E;    16'd52882: out <= 16'h0306;    16'd52883: out <= 16'h0291;
    16'd52884: out <= 16'h0272;    16'd52885: out <= 16'h017C;    16'd52886: out <= 16'h08F7;    16'd52887: out <= 16'h0031;
    16'd52888: out <= 16'h04EA;    16'd52889: out <= 16'h0399;    16'd52890: out <= 16'h047C;    16'd52891: out <= 16'h04DC;
    16'd52892: out <= 16'h04C5;    16'd52893: out <= 16'h0785;    16'd52894: out <= 16'h027C;    16'd52895: out <= 16'h05BB;
    16'd52896: out <= 16'h02D1;    16'd52897: out <= 16'h065F;    16'd52898: out <= 16'h0360;    16'd52899: out <= 16'h03D6;
    16'd52900: out <= 16'h00DC;    16'd52901: out <= 16'h0586;    16'd52902: out <= 16'h03B3;    16'd52903: out <= 16'h08B2;
    16'd52904: out <= 16'h09ED;    16'd52905: out <= 16'h0771;    16'd52906: out <= 16'h0069;    16'd52907: out <= 16'h01C5;
    16'd52908: out <= 16'h0ACD;    16'd52909: out <= 16'h090F;    16'd52910: out <= 16'h00B1;    16'd52911: out <= 16'h02D0;
    16'd52912: out <= 16'h028A;    16'd52913: out <= 16'h02C6;    16'd52914: out <= 16'h0153;    16'd52915: out <= 16'h05DA;
    16'd52916: out <= 16'h0926;    16'd52917: out <= 16'h027A;    16'd52918: out <= 16'h01A2;    16'd52919: out <= 16'hFF99;
    16'd52920: out <= 16'h02A9;    16'd52921: out <= 16'h0198;    16'd52922: out <= 16'h03D9;    16'd52923: out <= 16'h0692;
    16'd52924: out <= 16'h05BA;    16'd52925: out <= 16'h045B;    16'd52926: out <= 16'h031F;    16'd52927: out <= 16'h00F7;
    16'd52928: out <= 16'hFFF3;    16'd52929: out <= 16'h0269;    16'd52930: out <= 16'h0092;    16'd52931: out <= 16'hFEAE;
    16'd52932: out <= 16'h0301;    16'd52933: out <= 16'hFD95;    16'd52934: out <= 16'hFE79;    16'd52935: out <= 16'hF8D5;
    16'd52936: out <= 16'hFCDD;    16'd52937: out <= 16'h0517;    16'd52938: out <= 16'hF874;    16'd52939: out <= 16'h0284;
    16'd52940: out <= 16'hFA2A;    16'd52941: out <= 16'hFC5D;    16'd52942: out <= 16'hFAB9;    16'd52943: out <= 16'hFE90;
    16'd52944: out <= 16'h07B8;    16'd52945: out <= 16'hFF44;    16'd52946: out <= 16'hFE27;    16'd52947: out <= 16'hF8EA;
    16'd52948: out <= 16'h02D0;    16'd52949: out <= 16'h0044;    16'd52950: out <= 16'hFD45;    16'd52951: out <= 16'hFC5A;
    16'd52952: out <= 16'hFA1C;    16'd52953: out <= 16'h030F;    16'd52954: out <= 16'hF745;    16'd52955: out <= 16'h08A1;
    16'd52956: out <= 16'hFABA;    16'd52957: out <= 16'hFB04;    16'd52958: out <= 16'h0812;    16'd52959: out <= 16'h0516;
    16'd52960: out <= 16'hFAE4;    16'd52961: out <= 16'h02D1;    16'd52962: out <= 16'hFC1F;    16'd52963: out <= 16'h06E3;
    16'd52964: out <= 16'h01A5;    16'd52965: out <= 16'h0512;    16'd52966: out <= 16'hFFC5;    16'd52967: out <= 16'hFF22;
    16'd52968: out <= 16'h004B;    16'd52969: out <= 16'hFACA;    16'd52970: out <= 16'h039D;    16'd52971: out <= 16'h068F;
    16'd52972: out <= 16'hFD09;    16'd52973: out <= 16'hFD7D;    16'd52974: out <= 16'hFB99;    16'd52975: out <= 16'hFDB5;
    16'd52976: out <= 16'h01C4;    16'd52977: out <= 16'hFF52;    16'd52978: out <= 16'hFB32;    16'd52979: out <= 16'hFDF9;
    16'd52980: out <= 16'h033A;    16'd52981: out <= 16'h05DC;    16'd52982: out <= 16'h0257;    16'd52983: out <= 16'h0AF4;
    16'd52984: out <= 16'hF85B;    16'd52985: out <= 16'hFEDC;    16'd52986: out <= 16'h00D6;    16'd52987: out <= 16'hFF6D;
    16'd52988: out <= 16'h0666;    16'd52989: out <= 16'h02BE;    16'd52990: out <= 16'h01BB;    16'd52991: out <= 16'h0728;
    16'd52992: out <= 16'hFB8D;    16'd52993: out <= 16'h010B;    16'd52994: out <= 16'hFD3E;    16'd52995: out <= 16'hFE71;
    16'd52996: out <= 16'h01E0;    16'd52997: out <= 16'h02A3;    16'd52998: out <= 16'h034F;    16'd52999: out <= 16'h019A;
    16'd53000: out <= 16'hF5F8;    16'd53001: out <= 16'hFDE5;    16'd53002: out <= 16'h0183;    16'd53003: out <= 16'h01A4;
    16'd53004: out <= 16'hF88B;    16'd53005: out <= 16'hFB77;    16'd53006: out <= 16'h0561;    16'd53007: out <= 16'h02AF;
    16'd53008: out <= 16'hFCC2;    16'd53009: out <= 16'h0275;    16'd53010: out <= 16'hFF12;    16'd53011: out <= 16'h05FB;
    16'd53012: out <= 16'h03B9;    16'd53013: out <= 16'hFF7A;    16'd53014: out <= 16'h050E;    16'd53015: out <= 16'h0534;
    16'd53016: out <= 16'hFC65;    16'd53017: out <= 16'h04EB;    16'd53018: out <= 16'hFF1E;    16'd53019: out <= 16'h01C4;
    16'd53020: out <= 16'h0284;    16'd53021: out <= 16'hFEFF;    16'd53022: out <= 16'h000D;    16'd53023: out <= 16'hFD5F;
    16'd53024: out <= 16'hFEA8;    16'd53025: out <= 16'hFB0D;    16'd53026: out <= 16'hFFEB;    16'd53027: out <= 16'h0093;
    16'd53028: out <= 16'h0672;    16'd53029: out <= 16'hFEDE;    16'd53030: out <= 16'h01E8;    16'd53031: out <= 16'hFAD5;
    16'd53032: out <= 16'hF7E0;    16'd53033: out <= 16'hFAD4;    16'd53034: out <= 16'h0AD0;    16'd53035: out <= 16'hFDE6;
    16'd53036: out <= 16'h005C;    16'd53037: out <= 16'h0373;    16'd53038: out <= 16'h0AF3;    16'd53039: out <= 16'hFF38;
    16'd53040: out <= 16'h004F;    16'd53041: out <= 16'h06F4;    16'd53042: out <= 16'h068E;    16'd53043: out <= 16'h020A;
    16'd53044: out <= 16'h01F3;    16'd53045: out <= 16'h032C;    16'd53046: out <= 16'h0EA8;    16'd53047: out <= 16'hFD3C;
    16'd53048: out <= 16'h01EC;    16'd53049: out <= 16'h04E7;    16'd53050: out <= 16'h01AE;    16'd53051: out <= 16'h0B09;
    16'd53052: out <= 16'hFF30;    16'd53053: out <= 16'h010D;    16'd53054: out <= 16'h0588;    16'd53055: out <= 16'h00F4;
    16'd53056: out <= 16'h0108;    16'd53057: out <= 16'h0680;    16'd53058: out <= 16'h04B3;    16'd53059: out <= 16'h0216;
    16'd53060: out <= 16'h007C;    16'd53061: out <= 16'h0098;    16'd53062: out <= 16'h037B;    16'd53063: out <= 16'h0A0D;
    16'd53064: out <= 16'h04F3;    16'd53065: out <= 16'h081F;    16'd53066: out <= 16'h01C7;    16'd53067: out <= 16'h06FA;
    16'd53068: out <= 16'hFFA6;    16'd53069: out <= 16'h0406;    16'd53070: out <= 16'hFE04;    16'd53071: out <= 16'h00A7;
    16'd53072: out <= 16'h078E;    16'd53073: out <= 16'h00AD;    16'd53074: out <= 16'h03A2;    16'd53075: out <= 16'h01C6;
    16'd53076: out <= 16'h02D0;    16'd53077: out <= 16'h0435;    16'd53078: out <= 16'h0309;    16'd53079: out <= 16'hFE7F;
    16'd53080: out <= 16'h00D5;    16'd53081: out <= 16'h05D0;    16'd53082: out <= 16'h0C63;    16'd53083: out <= 16'h00CF;
    16'd53084: out <= 16'h0541;    16'd53085: out <= 16'hFD9A;    16'd53086: out <= 16'h01F7;    16'd53087: out <= 16'h06E5;
    16'd53088: out <= 16'hFE21;    16'd53089: out <= 16'hFCB2;    16'd53090: out <= 16'hFD8C;    16'd53091: out <= 16'hFFE4;
    16'd53092: out <= 16'h00BA;    16'd53093: out <= 16'h042C;    16'd53094: out <= 16'hFA3F;    16'd53095: out <= 16'h006D;
    16'd53096: out <= 16'h046C;    16'd53097: out <= 16'hFC5C;    16'd53098: out <= 16'h043F;    16'd53099: out <= 16'hFE7C;
    16'd53100: out <= 16'h0105;    16'd53101: out <= 16'hF61E;    16'd53102: out <= 16'h01C7;    16'd53103: out <= 16'hF8BF;
    16'd53104: out <= 16'hFE54;    16'd53105: out <= 16'hFCDE;    16'd53106: out <= 16'h024E;    16'd53107: out <= 16'h045D;
    16'd53108: out <= 16'h0292;    16'd53109: out <= 16'hFFC4;    16'd53110: out <= 16'hFDC3;    16'd53111: out <= 16'hFEFF;
    16'd53112: out <= 16'hFF37;    16'd53113: out <= 16'hFFAA;    16'd53114: out <= 16'h04E8;    16'd53115: out <= 16'h0198;
    16'd53116: out <= 16'hF8AB;    16'd53117: out <= 16'h0230;    16'd53118: out <= 16'h0D7D;    16'd53119: out <= 16'hFC0B;
    16'd53120: out <= 16'hFF3F;    16'd53121: out <= 16'hFC24;    16'd53122: out <= 16'h02B9;    16'd53123: out <= 16'h00A7;
    16'd53124: out <= 16'h093D;    16'd53125: out <= 16'h01DE;    16'd53126: out <= 16'h0586;    16'd53127: out <= 16'h03FD;
    16'd53128: out <= 16'h043E;    16'd53129: out <= 16'h02D1;    16'd53130: out <= 16'h08A2;    16'd53131: out <= 16'h011B;
    16'd53132: out <= 16'h04B4;    16'd53133: out <= 16'h0399;    16'd53134: out <= 16'h0A9A;    16'd53135: out <= 16'h008D;
    16'd53136: out <= 16'h0981;    16'd53137: out <= 16'h0846;    16'd53138: out <= 16'h0874;    16'd53139: out <= 16'h01FD;
    16'd53140: out <= 16'h0727;    16'd53141: out <= 16'h03D7;    16'd53142: out <= 16'h0682;    16'd53143: out <= 16'hFF3B;
    16'd53144: out <= 16'h025B;    16'd53145: out <= 16'h0024;    16'd53146: out <= 16'h08F2;    16'd53147: out <= 16'h031B;
    16'd53148: out <= 16'h091D;    16'd53149: out <= 16'hFEA2;    16'd53150: out <= 16'h02F4;    16'd53151: out <= 16'hFFBD;
    16'd53152: out <= 16'h0195;    16'd53153: out <= 16'h0675;    16'd53154: out <= 16'h031D;    16'd53155: out <= 16'hFA31;
    16'd53156: out <= 16'h0967;    16'd53157: out <= 16'h0105;    16'd53158: out <= 16'h02F9;    16'd53159: out <= 16'h0A83;
    16'd53160: out <= 16'h0177;    16'd53161: out <= 16'h091A;    16'd53162: out <= 16'h091E;    16'd53163: out <= 16'hFFDC;
    16'd53164: out <= 16'h092C;    16'd53165: out <= 16'h0268;    16'd53166: out <= 16'h09A8;    16'd53167: out <= 16'h009E;
    16'd53168: out <= 16'h055E;    16'd53169: out <= 16'h03FE;    16'd53170: out <= 16'h09A3;    16'd53171: out <= 16'h0054;
    16'd53172: out <= 16'h0365;    16'd53173: out <= 16'hFF9B;    16'd53174: out <= 16'h0345;    16'd53175: out <= 16'h0042;
    16'd53176: out <= 16'h02E3;    16'd53177: out <= 16'hFEAF;    16'd53178: out <= 16'h0550;    16'd53179: out <= 16'h0512;
    16'd53180: out <= 16'h0A58;    16'd53181: out <= 16'hFFDA;    16'd53182: out <= 16'h0497;    16'd53183: out <= 16'h069F;
    16'd53184: out <= 16'h0455;    16'd53185: out <= 16'h0664;    16'd53186: out <= 16'h0231;    16'd53187: out <= 16'h068F;
    16'd53188: out <= 16'h01C8;    16'd53189: out <= 16'hFBB0;    16'd53190: out <= 16'hFA8F;    16'd53191: out <= 16'hFC1A;
    16'd53192: out <= 16'hFFC5;    16'd53193: out <= 16'hF9A1;    16'd53194: out <= 16'hF849;    16'd53195: out <= 16'h0634;
    16'd53196: out <= 16'h0268;    16'd53197: out <= 16'h0443;    16'd53198: out <= 16'hFB2E;    16'd53199: out <= 16'h0340;
    16'd53200: out <= 16'h007B;    16'd53201: out <= 16'hFB73;    16'd53202: out <= 16'h0032;    16'd53203: out <= 16'h0494;
    16'd53204: out <= 16'hFE6C;    16'd53205: out <= 16'h017E;    16'd53206: out <= 16'hF8A5;    16'd53207: out <= 16'hFD26;
    16'd53208: out <= 16'h0303;    16'd53209: out <= 16'h0122;    16'd53210: out <= 16'hFD51;    16'd53211: out <= 16'hFF11;
    16'd53212: out <= 16'hFF36;    16'd53213: out <= 16'hFDFC;    16'd53214: out <= 16'hFE26;    16'd53215: out <= 16'hFC1D;
    16'd53216: out <= 16'hFEAF;    16'd53217: out <= 16'h02E5;    16'd53218: out <= 16'h0055;    16'd53219: out <= 16'h0753;
    16'd53220: out <= 16'hFF86;    16'd53221: out <= 16'hFDC9;    16'd53222: out <= 16'hFE3B;    16'd53223: out <= 16'hFCC8;
    16'd53224: out <= 16'h018A;    16'd53225: out <= 16'hFDBF;    16'd53226: out <= 16'h0083;    16'd53227: out <= 16'hF957;
    16'd53228: out <= 16'hFC8E;    16'd53229: out <= 16'h011D;    16'd53230: out <= 16'hFCEF;    16'd53231: out <= 16'hFCE6;
    16'd53232: out <= 16'h0100;    16'd53233: out <= 16'h0327;    16'd53234: out <= 16'hFC6C;    16'd53235: out <= 16'h0831;
    16'd53236: out <= 16'hFA8D;    16'd53237: out <= 16'hFE4B;    16'd53238: out <= 16'hFA3E;    16'd53239: out <= 16'hFD6B;
    16'd53240: out <= 16'hFE5A;    16'd53241: out <= 16'hFF9E;    16'd53242: out <= 16'h0001;    16'd53243: out <= 16'hF9A4;
    16'd53244: out <= 16'hFB14;    16'd53245: out <= 16'hFF49;    16'd53246: out <= 16'h0359;    16'd53247: out <= 16'hFCC5;
    16'd53248: out <= 16'hFC3A;    16'd53249: out <= 16'h0134;    16'd53250: out <= 16'h027E;    16'd53251: out <= 16'hFC3B;
    16'd53252: out <= 16'hFF2B;    16'd53253: out <= 16'hFFCD;    16'd53254: out <= 16'h063C;    16'd53255: out <= 16'hFC33;
    16'd53256: out <= 16'hFA7F;    16'd53257: out <= 16'h02B8;    16'd53258: out <= 16'h06BD;    16'd53259: out <= 16'h0272;
    16'd53260: out <= 16'hFFF1;    16'd53261: out <= 16'h0484;    16'd53262: out <= 16'h0B19;    16'd53263: out <= 16'h053B;
    16'd53264: out <= 16'h0088;    16'd53265: out <= 16'h0327;    16'd53266: out <= 16'h0746;    16'd53267: out <= 16'hFB44;
    16'd53268: out <= 16'h038A;    16'd53269: out <= 16'hFD35;    16'd53270: out <= 16'hF965;    16'd53271: out <= 16'h008E;
    16'd53272: out <= 16'h044B;    16'd53273: out <= 16'hFCE2;    16'd53274: out <= 16'h00AF;    16'd53275: out <= 16'h0194;
    16'd53276: out <= 16'hFD60;    16'd53277: out <= 16'h06E1;    16'd53278: out <= 16'h056C;    16'd53279: out <= 16'h02DF;
    16'd53280: out <= 16'h044E;    16'd53281: out <= 16'hFEB2;    16'd53282: out <= 16'hFEE4;    16'd53283: out <= 16'h0346;
    16'd53284: out <= 16'h03CC;    16'd53285: out <= 16'h026A;    16'd53286: out <= 16'h075E;    16'd53287: out <= 16'hFEEE;
    16'd53288: out <= 16'hF745;    16'd53289: out <= 16'h0315;    16'd53290: out <= 16'hFD55;    16'd53291: out <= 16'h0446;
    16'd53292: out <= 16'h01AA;    16'd53293: out <= 16'h017F;    16'd53294: out <= 16'hFDB0;    16'd53295: out <= 16'hFE23;
    16'd53296: out <= 16'h0AE9;    16'd53297: out <= 16'h099F;    16'd53298: out <= 16'hFD76;    16'd53299: out <= 16'h0175;
    16'd53300: out <= 16'h0078;    16'd53301: out <= 16'h02D4;    16'd53302: out <= 16'h0121;    16'd53303: out <= 16'h0B5C;
    16'd53304: out <= 16'h07B6;    16'd53305: out <= 16'hFF76;    16'd53306: out <= 16'h0277;    16'd53307: out <= 16'h0355;
    16'd53308: out <= 16'h00B3;    16'd53309: out <= 16'h004E;    16'd53310: out <= 16'h0878;    16'd53311: out <= 16'h04FA;
    16'd53312: out <= 16'h0791;    16'd53313: out <= 16'h0168;    16'd53314: out <= 16'h01E7;    16'd53315: out <= 16'hFE89;
    16'd53316: out <= 16'h0A7B;    16'd53317: out <= 16'h0621;    16'd53318: out <= 16'hFF8E;    16'd53319: out <= 16'h0308;
    16'd53320: out <= 16'h01C2;    16'd53321: out <= 16'h0E1D;    16'd53322: out <= 16'h0540;    16'd53323: out <= 16'h004F;
    16'd53324: out <= 16'h0465;    16'd53325: out <= 16'hFF0F;    16'd53326: out <= 16'h0498;    16'd53327: out <= 16'h03A0;
    16'd53328: out <= 16'h0288;    16'd53329: out <= 16'h0343;    16'd53330: out <= 16'h04C5;    16'd53331: out <= 16'h03A7;
    16'd53332: out <= 16'h0438;    16'd53333: out <= 16'h0461;    16'd53334: out <= 16'h0998;    16'd53335: out <= 16'h0547;
    16'd53336: out <= 16'h059D;    16'd53337: out <= 16'h0C17;    16'd53338: out <= 16'h0757;    16'd53339: out <= 16'h02DD;
    16'd53340: out <= 16'hFD6D;    16'd53341: out <= 16'h030C;    16'd53342: out <= 16'h0AEB;    16'd53343: out <= 16'hFE14;
    16'd53344: out <= 16'hFEB0;    16'd53345: out <= 16'h0431;    16'd53346: out <= 16'h015E;    16'd53347: out <= 16'hFFBB;
    16'd53348: out <= 16'h03CD;    16'd53349: out <= 16'h0136;    16'd53350: out <= 16'hFB2A;    16'd53351: out <= 16'h0087;
    16'd53352: out <= 16'hFDB9;    16'd53353: out <= 16'h05BF;    16'd53354: out <= 16'hFF88;    16'd53355: out <= 16'hF944;
    16'd53356: out <= 16'hFF2B;    16'd53357: out <= 16'h0150;    16'd53358: out <= 16'h0102;    16'd53359: out <= 16'hFE6C;
    16'd53360: out <= 16'h060F;    16'd53361: out <= 16'hFDEA;    16'd53362: out <= 16'hFEA2;    16'd53363: out <= 16'h00D9;
    16'd53364: out <= 16'hFD17;    16'd53365: out <= 16'h04FE;    16'd53366: out <= 16'h03CA;    16'd53367: out <= 16'hFC70;
    16'd53368: out <= 16'h06F0;    16'd53369: out <= 16'h0223;    16'd53370: out <= 16'h01DD;    16'd53371: out <= 16'hFDAB;
    16'd53372: out <= 16'hFB47;    16'd53373: out <= 16'hFE4D;    16'd53374: out <= 16'h02A1;    16'd53375: out <= 16'hFF25;
    16'd53376: out <= 16'h00B0;    16'd53377: out <= 16'h024E;    16'd53378: out <= 16'hFBA4;    16'd53379: out <= 16'hFB73;
    16'd53380: out <= 16'h00FE;    16'd53381: out <= 16'h028B;    16'd53382: out <= 16'h0021;    16'd53383: out <= 16'hFC30;
    16'd53384: out <= 16'h01BD;    16'd53385: out <= 16'h0933;    16'd53386: out <= 16'h038C;    16'd53387: out <= 16'h02C0;
    16'd53388: out <= 16'h052A;    16'd53389: out <= 16'hFAC8;    16'd53390: out <= 16'h02FA;    16'd53391: out <= 16'h0A08;
    16'd53392: out <= 16'h05AE;    16'd53393: out <= 16'h0755;    16'd53394: out <= 16'h01DD;    16'd53395: out <= 16'h080F;
    16'd53396: out <= 16'h040B;    16'd53397: out <= 16'h04D6;    16'd53398: out <= 16'h01B3;    16'd53399: out <= 16'h01CB;
    16'd53400: out <= 16'h03F7;    16'd53401: out <= 16'h0906;    16'd53402: out <= 16'h0588;    16'd53403: out <= 16'h0E6D;
    16'd53404: out <= 16'h01D1;    16'd53405: out <= 16'h06FE;    16'd53406: out <= 16'h03CF;    16'd53407: out <= 16'hFED0;
    16'd53408: out <= 16'hFB04;    16'd53409: out <= 16'h0287;    16'd53410: out <= 16'h035C;    16'd53411: out <= 16'h01A8;
    16'd53412: out <= 16'h0048;    16'd53413: out <= 16'h01AA;    16'd53414: out <= 16'h05B1;    16'd53415: out <= 16'h034C;
    16'd53416: out <= 16'h023F;    16'd53417: out <= 16'h0396;    16'd53418: out <= 16'h0700;    16'd53419: out <= 16'h0165;
    16'd53420: out <= 16'h0818;    16'd53421: out <= 16'h0BAD;    16'd53422: out <= 16'h0063;    16'd53423: out <= 16'hFC5F;
    16'd53424: out <= 16'h0002;    16'd53425: out <= 16'h021E;    16'd53426: out <= 16'h0050;    16'd53427: out <= 16'h050A;
    16'd53428: out <= 16'h04EC;    16'd53429: out <= 16'h01AB;    16'd53430: out <= 16'hFC4E;    16'd53431: out <= 16'h0FFB;
    16'd53432: out <= 16'h020B;    16'd53433: out <= 16'h01F0;    16'd53434: out <= 16'hFE29;    16'd53435: out <= 16'h04AA;
    16'd53436: out <= 16'h078B;    16'd53437: out <= 16'h03FC;    16'd53438: out <= 16'hFF27;    16'd53439: out <= 16'h02AE;
    16'd53440: out <= 16'h023B;    16'd53441: out <= 16'h00B9;    16'd53442: out <= 16'h035E;    16'd53443: out <= 16'hF857;
    16'd53444: out <= 16'hFEC9;    16'd53445: out <= 16'h0380;    16'd53446: out <= 16'h001D;    16'd53447: out <= 16'hFE64;
    16'd53448: out <= 16'hFFF6;    16'd53449: out <= 16'hFF30;    16'd53450: out <= 16'h0B10;    16'd53451: out <= 16'h036B;
    16'd53452: out <= 16'hFD47;    16'd53453: out <= 16'h0321;    16'd53454: out <= 16'h08E3;    16'd53455: out <= 16'h005E;
    16'd53456: out <= 16'h000A;    16'd53457: out <= 16'hFCCD;    16'd53458: out <= 16'h02A8;    16'd53459: out <= 16'hFC6F;
    16'd53460: out <= 16'h05A2;    16'd53461: out <= 16'h0214;    16'd53462: out <= 16'hF991;    16'd53463: out <= 16'hFF80;
    16'd53464: out <= 16'h0192;    16'd53465: out <= 16'h04BF;    16'd53466: out <= 16'h0453;    16'd53467: out <= 16'hFF29;
    16'd53468: out <= 16'hFB95;    16'd53469: out <= 16'hFA22;    16'd53470: out <= 16'h01E0;    16'd53471: out <= 16'h0397;
    16'd53472: out <= 16'hF9EB;    16'd53473: out <= 16'hFFE9;    16'd53474: out <= 16'h0802;    16'd53475: out <= 16'hFEE8;
    16'd53476: out <= 16'h00F9;    16'd53477: out <= 16'h053B;    16'd53478: out <= 16'hFEA6;    16'd53479: out <= 16'hFD2F;
    16'd53480: out <= 16'hF538;    16'd53481: out <= 16'hFF96;    16'd53482: out <= 16'hF62E;    16'd53483: out <= 16'h02DB;
    16'd53484: out <= 16'h02BE;    16'd53485: out <= 16'hFB81;    16'd53486: out <= 16'hFD87;    16'd53487: out <= 16'hFAF8;
    16'd53488: out <= 16'h01C7;    16'd53489: out <= 16'h04D7;    16'd53490: out <= 16'h0153;    16'd53491: out <= 16'hFC87;
    16'd53492: out <= 16'h026B;    16'd53493: out <= 16'hFE01;    16'd53494: out <= 16'hFA05;    16'd53495: out <= 16'h0547;
    16'd53496: out <= 16'hF73B;    16'd53497: out <= 16'h03D9;    16'd53498: out <= 16'h0007;    16'd53499: out <= 16'h012D;
    16'd53500: out <= 16'h039A;    16'd53501: out <= 16'h054E;    16'd53502: out <= 16'h0088;    16'd53503: out <= 16'hFE5F;
    16'd53504: out <= 16'h0150;    16'd53505: out <= 16'h011E;    16'd53506: out <= 16'h00CE;    16'd53507: out <= 16'hFA1D;
    16'd53508: out <= 16'h0072;    16'd53509: out <= 16'hFFEA;    16'd53510: out <= 16'hF79A;    16'd53511: out <= 16'hFFAC;
    16'd53512: out <= 16'hF9D9;    16'd53513: out <= 16'h01A4;    16'd53514: out <= 16'h02D3;    16'd53515: out <= 16'hFFA9;
    16'd53516: out <= 16'h019E;    16'd53517: out <= 16'h01DF;    16'd53518: out <= 16'h018C;    16'd53519: out <= 16'hF836;
    16'd53520: out <= 16'h0582;    16'd53521: out <= 16'hFA4C;    16'd53522: out <= 16'hFD94;    16'd53523: out <= 16'hFF92;
    16'd53524: out <= 16'h00F0;    16'd53525: out <= 16'hFF90;    16'd53526: out <= 16'hFBF4;    16'd53527: out <= 16'h027F;
    16'd53528: out <= 16'h0352;    16'd53529: out <= 16'h02B9;    16'd53530: out <= 16'h0044;    16'd53531: out <= 16'hFE2C;
    16'd53532: out <= 16'hFF92;    16'd53533: out <= 16'h0352;    16'd53534: out <= 16'hFFF0;    16'd53535: out <= 16'hF8A3;
    16'd53536: out <= 16'hFF4F;    16'd53537: out <= 16'h0387;    16'd53538: out <= 16'hFCF0;    16'd53539: out <= 16'hFD17;
    16'd53540: out <= 16'h056F;    16'd53541: out <= 16'hFC90;    16'd53542: out <= 16'hFF9A;    16'd53543: out <= 16'hFE0B;
    16'd53544: out <= 16'h063E;    16'd53545: out <= 16'h062F;    16'd53546: out <= 16'h064C;    16'd53547: out <= 16'h0229;
    16'd53548: out <= 16'hFA0C;    16'd53549: out <= 16'h077F;    16'd53550: out <= 16'hFABC;    16'd53551: out <= 16'hF829;
    16'd53552: out <= 16'hFD82;    16'd53553: out <= 16'h0588;    16'd53554: out <= 16'h0156;    16'd53555: out <= 16'h0551;
    16'd53556: out <= 16'h0166;    16'd53557: out <= 16'h06EB;    16'd53558: out <= 16'h0769;    16'd53559: out <= 16'h07BB;
    16'd53560: out <= 16'h0561;    16'd53561: out <= 16'h07CA;    16'd53562: out <= 16'h0263;    16'd53563: out <= 16'h0100;
    16'd53564: out <= 16'h0A20;    16'd53565: out <= 16'h0018;    16'd53566: out <= 16'hFA1E;    16'd53567: out <= 16'h038E;
    16'd53568: out <= 16'hFE53;    16'd53569: out <= 16'h0165;    16'd53570: out <= 16'h01ED;    16'd53571: out <= 16'h0396;
    16'd53572: out <= 16'h071B;    16'd53573: out <= 16'h0639;    16'd53574: out <= 16'h047D;    16'd53575: out <= 16'h00AE;
    16'd53576: out <= 16'h07DA;    16'd53577: out <= 16'h0891;    16'd53578: out <= 16'h05FC;    16'd53579: out <= 16'h0598;
    16'd53580: out <= 16'hFC9A;    16'd53581: out <= 16'h06D4;    16'd53582: out <= 16'hFD97;    16'd53583: out <= 16'h06D1;
    16'd53584: out <= 16'h0563;    16'd53585: out <= 16'h037D;    16'd53586: out <= 16'hFA83;    16'd53587: out <= 16'h0762;
    16'd53588: out <= 16'h03DA;    16'd53589: out <= 16'h033E;    16'd53590: out <= 16'h05A8;    16'd53591: out <= 16'h068E;
    16'd53592: out <= 16'h02F5;    16'd53593: out <= 16'h0663;    16'd53594: out <= 16'h03A9;    16'd53595: out <= 16'hFE10;
    16'd53596: out <= 16'hFE4E;    16'd53597: out <= 16'hFC98;    16'd53598: out <= 16'h06E9;    16'd53599: out <= 16'h0133;
    16'd53600: out <= 16'hFD67;    16'd53601: out <= 16'hFE4B;    16'd53602: out <= 16'hFFB7;    16'd53603: out <= 16'hF843;
    16'd53604: out <= 16'hFB17;    16'd53605: out <= 16'hFE5E;    16'd53606: out <= 16'h0131;    16'd53607: out <= 16'hFD5B;
    16'd53608: out <= 16'h04CA;    16'd53609: out <= 16'h0379;    16'd53610: out <= 16'h005E;    16'd53611: out <= 16'hFFC3;
    16'd53612: out <= 16'hFBFA;    16'd53613: out <= 16'hFF64;    16'd53614: out <= 16'h0436;    16'd53615: out <= 16'hFE9D;
    16'd53616: out <= 16'hFA90;    16'd53617: out <= 16'hFBB9;    16'd53618: out <= 16'hFFED;    16'd53619: out <= 16'hF901;
    16'd53620: out <= 16'h044D;    16'd53621: out <= 16'h0064;    16'd53622: out <= 16'hFA84;    16'd53623: out <= 16'hFF8C;
    16'd53624: out <= 16'hFE29;    16'd53625: out <= 16'h01E2;    16'd53626: out <= 16'h0531;    16'd53627: out <= 16'h009E;
    16'd53628: out <= 16'h00BB;    16'd53629: out <= 16'hFE8B;    16'd53630: out <= 16'h035B;    16'd53631: out <= 16'hFD1F;
    16'd53632: out <= 16'hFCD2;    16'd53633: out <= 16'hFCF9;    16'd53634: out <= 16'hFD95;    16'd53635: out <= 16'h018C;
    16'd53636: out <= 16'h084D;    16'd53637: out <= 16'h0709;    16'd53638: out <= 16'h008A;    16'd53639: out <= 16'hFF46;
    16'd53640: out <= 16'hFE7A;    16'd53641: out <= 16'h00A0;    16'd53642: out <= 16'h0242;    16'd53643: out <= 16'hFFBB;
    16'd53644: out <= 16'h02BA;    16'd53645: out <= 16'h06D0;    16'd53646: out <= 16'h0548;    16'd53647: out <= 16'h04F3;
    16'd53648: out <= 16'h01A5;    16'd53649: out <= 16'h090F;    16'd53650: out <= 16'h0609;    16'd53651: out <= 16'hFFB0;
    16'd53652: out <= 16'h0AF2;    16'd53653: out <= 16'hFDEC;    16'd53654: out <= 16'hFF49;    16'd53655: out <= 16'hFF67;
    16'd53656: out <= 16'h0168;    16'd53657: out <= 16'h0336;    16'd53658: out <= 16'h06F3;    16'd53659: out <= 16'h07F1;
    16'd53660: out <= 16'h07E6;    16'd53661: out <= 16'h04E4;    16'd53662: out <= 16'h08CA;    16'd53663: out <= 16'h0024;
    16'd53664: out <= 16'h00DE;    16'd53665: out <= 16'h029A;    16'd53666: out <= 16'h0443;    16'd53667: out <= 16'hFED1;
    16'd53668: out <= 16'h0573;    16'd53669: out <= 16'hFB24;    16'd53670: out <= 16'h023D;    16'd53671: out <= 16'hFE0A;
    16'd53672: out <= 16'hFEBF;    16'd53673: out <= 16'h070F;    16'd53674: out <= 16'h09DB;    16'd53675: out <= 16'h0972;
    16'd53676: out <= 16'h04D5;    16'd53677: out <= 16'h041E;    16'd53678: out <= 16'h023F;    16'd53679: out <= 16'hFA83;
    16'd53680: out <= 16'h0313;    16'd53681: out <= 16'h0150;    16'd53682: out <= 16'h02CC;    16'd53683: out <= 16'h09EF;
    16'd53684: out <= 16'h07A5;    16'd53685: out <= 16'h0717;    16'd53686: out <= 16'h0985;    16'd53687: out <= 16'h0423;
    16'd53688: out <= 16'h01D4;    16'd53689: out <= 16'h01D5;    16'd53690: out <= 16'h0C2C;    16'd53691: out <= 16'h0887;
    16'd53692: out <= 16'h0584;    16'd53693: out <= 16'h0394;    16'd53694: out <= 16'h000A;    16'd53695: out <= 16'h04A0;
    16'd53696: out <= 16'h0454;    16'd53697: out <= 16'h08A2;    16'd53698: out <= 16'h03A7;    16'd53699: out <= 16'h02FD;
    16'd53700: out <= 16'h045E;    16'd53701: out <= 16'h03A5;    16'd53702: out <= 16'h0069;    16'd53703: out <= 16'h03EE;
    16'd53704: out <= 16'hFC1F;    16'd53705: out <= 16'h041C;    16'd53706: out <= 16'h0455;    16'd53707: out <= 16'h03E6;
    16'd53708: out <= 16'h048A;    16'd53709: out <= 16'h0201;    16'd53710: out <= 16'hFCFE;    16'd53711: out <= 16'hFC5F;
    16'd53712: out <= 16'h0077;    16'd53713: out <= 16'h0297;    16'd53714: out <= 16'hFE82;    16'd53715: out <= 16'h055E;
    16'd53716: out <= 16'hFE7D;    16'd53717: out <= 16'h0125;    16'd53718: out <= 16'h01F2;    16'd53719: out <= 16'hFF18;
    16'd53720: out <= 16'hFD3C;    16'd53721: out <= 16'h0246;    16'd53722: out <= 16'h0348;    16'd53723: out <= 16'hFF4A;
    16'd53724: out <= 16'h0140;    16'd53725: out <= 16'hFD41;    16'd53726: out <= 16'hFEC3;    16'd53727: out <= 16'hFC90;
    16'd53728: out <= 16'h0280;    16'd53729: out <= 16'hFFDF;    16'd53730: out <= 16'hFACE;    16'd53731: out <= 16'hFDDE;
    16'd53732: out <= 16'hF87B;    16'd53733: out <= 16'hFB6E;    16'd53734: out <= 16'h0461;    16'd53735: out <= 16'hF91C;
    16'd53736: out <= 16'hFD65;    16'd53737: out <= 16'hFF89;    16'd53738: out <= 16'h083C;    16'd53739: out <= 16'hFE72;
    16'd53740: out <= 16'hFF67;    16'd53741: out <= 16'h0211;    16'd53742: out <= 16'h0690;    16'd53743: out <= 16'h014F;
    16'd53744: out <= 16'h03F6;    16'd53745: out <= 16'hFC44;    16'd53746: out <= 16'h0366;    16'd53747: out <= 16'hFF6C;
    16'd53748: out <= 16'hFF8A;    16'd53749: out <= 16'h0479;    16'd53750: out <= 16'h0061;    16'd53751: out <= 16'hFEDE;
    16'd53752: out <= 16'hFCD4;    16'd53753: out <= 16'h018F;    16'd53754: out <= 16'hF711;    16'd53755: out <= 16'h09F8;
    16'd53756: out <= 16'h0336;    16'd53757: out <= 16'h016C;    16'd53758: out <= 16'h016F;    16'd53759: out <= 16'hFFB1;
    16'd53760: out <= 16'h0525;    16'd53761: out <= 16'hFE0A;    16'd53762: out <= 16'hFC47;    16'd53763: out <= 16'h007E;
    16'd53764: out <= 16'h037E;    16'd53765: out <= 16'hF76E;    16'd53766: out <= 16'hFF80;    16'd53767: out <= 16'h080D;
    16'd53768: out <= 16'hFEF3;    16'd53769: out <= 16'h02DD;    16'd53770: out <= 16'h03E0;    16'd53771: out <= 16'h0447;
    16'd53772: out <= 16'hFECC;    16'd53773: out <= 16'hFB48;    16'd53774: out <= 16'hFE6A;    16'd53775: out <= 16'hFE6F;
    16'd53776: out <= 16'hFE20;    16'd53777: out <= 16'h0525;    16'd53778: out <= 16'hFE8A;    16'd53779: out <= 16'h0056;
    16'd53780: out <= 16'hFE1A;    16'd53781: out <= 16'h00F7;    16'd53782: out <= 16'hF84D;    16'd53783: out <= 16'h031B;
    16'd53784: out <= 16'h02E2;    16'd53785: out <= 16'h07B3;    16'd53786: out <= 16'h05BA;    16'd53787: out <= 16'hFD9F;
    16'd53788: out <= 16'hFE94;    16'd53789: out <= 16'hFA3F;    16'd53790: out <= 16'h04D7;    16'd53791: out <= 16'h03AC;
    16'd53792: out <= 16'hFBFF;    16'd53793: out <= 16'h03CA;    16'd53794: out <= 16'h0443;    16'd53795: out <= 16'hFA1F;
    16'd53796: out <= 16'hFE63;    16'd53797: out <= 16'hFDEB;    16'd53798: out <= 16'h0108;    16'd53799: out <= 16'h039E;
    16'd53800: out <= 16'hFB99;    16'd53801: out <= 16'hFF46;    16'd53802: out <= 16'hFD7D;    16'd53803: out <= 16'h00D3;
    16'd53804: out <= 16'h001F;    16'd53805: out <= 16'hFD28;    16'd53806: out <= 16'h0245;    16'd53807: out <= 16'h03C9;
    16'd53808: out <= 16'h049E;    16'd53809: out <= 16'hFF5C;    16'd53810: out <= 16'h0505;    16'd53811: out <= 16'h0599;
    16'd53812: out <= 16'h0A4D;    16'd53813: out <= 16'h06C7;    16'd53814: out <= 16'hFF19;    16'd53815: out <= 16'h03F2;
    16'd53816: out <= 16'hFCE4;    16'd53817: out <= 16'hFC2C;    16'd53818: out <= 16'h0B7B;    16'd53819: out <= 16'h026A;
    16'd53820: out <= 16'hF9A0;    16'd53821: out <= 16'h039F;    16'd53822: out <= 16'h039A;    16'd53823: out <= 16'h0004;
    16'd53824: out <= 16'h038D;    16'd53825: out <= 16'h032B;    16'd53826: out <= 16'hFFC0;    16'd53827: out <= 16'hFEE3;
    16'd53828: out <= 16'h07C3;    16'd53829: out <= 16'h03D0;    16'd53830: out <= 16'h01A2;    16'd53831: out <= 16'h02B6;
    16'd53832: out <= 16'h052B;    16'd53833: out <= 16'h0477;    16'd53834: out <= 16'h039A;    16'd53835: out <= 16'h0A66;
    16'd53836: out <= 16'h07A1;    16'd53837: out <= 16'h042A;    16'd53838: out <= 16'h0631;    16'd53839: out <= 16'hFC58;
    16'd53840: out <= 16'h01D8;    16'd53841: out <= 16'h032B;    16'd53842: out <= 16'hFCDA;    16'd53843: out <= 16'h0384;
    16'd53844: out <= 16'h0554;    16'd53845: out <= 16'h0625;    16'd53846: out <= 16'h0B29;    16'd53847: out <= 16'h044D;
    16'd53848: out <= 16'h0535;    16'd53849: out <= 16'h0182;    16'd53850: out <= 16'h07FD;    16'd53851: out <= 16'h0481;
    16'd53852: out <= 16'h06AD;    16'd53853: out <= 16'hFF7A;    16'd53854: out <= 16'h02AC;    16'd53855: out <= 16'h047D;
    16'd53856: out <= 16'h0156;    16'd53857: out <= 16'h01E4;    16'd53858: out <= 16'h0396;    16'd53859: out <= 16'hFF82;
    16'd53860: out <= 16'h02DD;    16'd53861: out <= 16'hF8A1;    16'd53862: out <= 16'hF83F;    16'd53863: out <= 16'hFF8C;
    16'd53864: out <= 16'hFD40;    16'd53865: out <= 16'h01E5;    16'd53866: out <= 16'h019E;    16'd53867: out <= 16'hFEC3;
    16'd53868: out <= 16'hF77B;    16'd53869: out <= 16'hF9D7;    16'd53870: out <= 16'h0567;    16'd53871: out <= 16'h02AC;
    16'd53872: out <= 16'h0257;    16'd53873: out <= 16'hFEE6;    16'd53874: out <= 16'h027D;    16'd53875: out <= 16'hFBE2;
    16'd53876: out <= 16'hFDD1;    16'd53877: out <= 16'h049F;    16'd53878: out <= 16'h00B7;    16'd53879: out <= 16'h0101;
    16'd53880: out <= 16'hFE69;    16'd53881: out <= 16'hFB7E;    16'd53882: out <= 16'h01A0;    16'd53883: out <= 16'hFD50;
    16'd53884: out <= 16'hFBA6;    16'd53885: out <= 16'h012A;    16'd53886: out <= 16'hFACE;    16'd53887: out <= 16'hFF74;
    16'd53888: out <= 16'hFF5B;    16'd53889: out <= 16'h01FB;    16'd53890: out <= 16'h057B;    16'd53891: out <= 16'h03FA;
    16'd53892: out <= 16'h025C;    16'd53893: out <= 16'h0011;    16'd53894: out <= 16'h0A55;    16'd53895: out <= 16'h0598;
    16'd53896: out <= 16'h04E9;    16'd53897: out <= 16'h00E5;    16'd53898: out <= 16'h0564;    16'd53899: out <= 16'h070E;
    16'd53900: out <= 16'h060E;    16'd53901: out <= 16'h09E8;    16'd53902: out <= 16'h0697;    16'd53903: out <= 16'h022F;
    16'd53904: out <= 16'h04B3;    16'd53905: out <= 16'h0734;    16'd53906: out <= 16'h001D;    16'd53907: out <= 16'h024C;
    16'd53908: out <= 16'h02FB;    16'd53909: out <= 16'h0657;    16'd53910: out <= 16'h031F;    16'd53911: out <= 16'h02BF;
    16'd53912: out <= 16'h00E6;    16'd53913: out <= 16'h056C;    16'd53914: out <= 16'h04ED;    16'd53915: out <= 16'h0396;
    16'd53916: out <= 16'h04F5;    16'd53917: out <= 16'h02B3;    16'd53918: out <= 16'h0A2E;    16'd53919: out <= 16'h0390;
    16'd53920: out <= 16'h0535;    16'd53921: out <= 16'hFCDD;    16'd53922: out <= 16'h05DC;    16'd53923: out <= 16'h08D7;
    16'd53924: out <= 16'h0081;    16'd53925: out <= 16'h017D;    16'd53926: out <= 16'h02EA;    16'd53927: out <= 16'h00C0;
    16'd53928: out <= 16'h0324;    16'd53929: out <= 16'h0333;    16'd53930: out <= 16'h0797;    16'd53931: out <= 16'h070F;
    16'd53932: out <= 16'h0658;    16'd53933: out <= 16'h02A7;    16'd53934: out <= 16'hFF9C;    16'd53935: out <= 16'h042E;
    16'd53936: out <= 16'h088B;    16'd53937: out <= 16'hFF98;    16'd53938: out <= 16'h0BAD;    16'd53939: out <= 16'h05B4;
    16'd53940: out <= 16'hFF98;    16'd53941: out <= 16'h06E7;    16'd53942: out <= 16'h041B;    16'd53943: out <= 16'h0245;
    16'd53944: out <= 16'h066B;    16'd53945: out <= 16'h0369;    16'd53946: out <= 16'h0AEB;    16'd53947: out <= 16'h05EC;
    16'd53948: out <= 16'h032A;    16'd53949: out <= 16'h0630;    16'd53950: out <= 16'h04EF;    16'd53951: out <= 16'h024C;
    16'd53952: out <= 16'h01F8;    16'd53953: out <= 16'hFED8;    16'd53954: out <= 16'h07DF;    16'd53955: out <= 16'hFF6B;
    16'd53956: out <= 16'hF6C7;    16'd53957: out <= 16'hFCEB;    16'd53958: out <= 16'hFB5E;    16'd53959: out <= 16'h0158;
    16'd53960: out <= 16'h0150;    16'd53961: out <= 16'h055D;    16'd53962: out <= 16'hFC86;    16'd53963: out <= 16'h0231;
    16'd53964: out <= 16'hFDBC;    16'd53965: out <= 16'hFDA2;    16'd53966: out <= 16'hF825;    16'd53967: out <= 16'h08C2;
    16'd53968: out <= 16'h031B;    16'd53969: out <= 16'h0322;    16'd53970: out <= 16'hFC69;    16'd53971: out <= 16'h053E;
    16'd53972: out <= 16'hFBED;    16'd53973: out <= 16'h033A;    16'd53974: out <= 16'hFC49;    16'd53975: out <= 16'h00DF;
    16'd53976: out <= 16'hFE21;    16'd53977: out <= 16'h00D7;    16'd53978: out <= 16'h01F6;    16'd53979: out <= 16'h0178;
    16'd53980: out <= 16'hF92B;    16'd53981: out <= 16'h031A;    16'd53982: out <= 16'hFF1C;    16'd53983: out <= 16'h011F;
    16'd53984: out <= 16'h0730;    16'd53985: out <= 16'hFF45;    16'd53986: out <= 16'hFBB7;    16'd53987: out <= 16'hFE08;
    16'd53988: out <= 16'h064E;    16'd53989: out <= 16'h003D;    16'd53990: out <= 16'hF91E;    16'd53991: out <= 16'hFB6B;
    16'd53992: out <= 16'hFCC2;    16'd53993: out <= 16'h00C3;    16'd53994: out <= 16'h025C;    16'd53995: out <= 16'hFFE9;
    16'd53996: out <= 16'h0173;    16'd53997: out <= 16'hFF3B;    16'd53998: out <= 16'h0185;    16'd53999: out <= 16'hFF1A;
    16'd54000: out <= 16'h0182;    16'd54001: out <= 16'hFAA4;    16'd54002: out <= 16'h0023;    16'd54003: out <= 16'hFD0E;
    16'd54004: out <= 16'hFFC5;    16'd54005: out <= 16'h06F2;    16'd54006: out <= 16'hF72A;    16'd54007: out <= 16'h02E8;
    16'd54008: out <= 16'h0179;    16'd54009: out <= 16'h032C;    16'd54010: out <= 16'hFE1A;    16'd54011: out <= 16'hFFC0;
    16'd54012: out <= 16'h0584;    16'd54013: out <= 16'hFED0;    16'd54014: out <= 16'h03C1;    16'd54015: out <= 16'hFFC2;
    16'd54016: out <= 16'hFED3;    16'd54017: out <= 16'h01ED;    16'd54018: out <= 16'hFE01;    16'd54019: out <= 16'hFE5C;
    16'd54020: out <= 16'hFDA7;    16'd54021: out <= 16'h029F;    16'd54022: out <= 16'h07A6;    16'd54023: out <= 16'hF8DF;
    16'd54024: out <= 16'h003C;    16'd54025: out <= 16'h0594;    16'd54026: out <= 16'hFD79;    16'd54027: out <= 16'hFDF6;
    16'd54028: out <= 16'h01DA;    16'd54029: out <= 16'hFB2F;    16'd54030: out <= 16'h02CD;    16'd54031: out <= 16'hFCD9;
    16'd54032: out <= 16'hFD4D;    16'd54033: out <= 16'h052B;    16'd54034: out <= 16'hFC58;    16'd54035: out <= 16'h0815;
    16'd54036: out <= 16'hFEE9;    16'd54037: out <= 16'hFCAC;    16'd54038: out <= 16'h00AE;    16'd54039: out <= 16'h05A4;
    16'd54040: out <= 16'h01FB;    16'd54041: out <= 16'h045A;    16'd54042: out <= 16'h012F;    16'd54043: out <= 16'h011D;
    16'd54044: out <= 16'h0289;    16'd54045: out <= 16'h00EC;    16'd54046: out <= 16'hFC23;    16'd54047: out <= 16'h03E7;
    16'd54048: out <= 16'h0538;    16'd54049: out <= 16'h04A6;    16'd54050: out <= 16'h095F;    16'd54051: out <= 16'hFF97;
    16'd54052: out <= 16'h065C;    16'd54053: out <= 16'hF879;    16'd54054: out <= 16'hFDE9;    16'd54055: out <= 16'hFA38;
    16'd54056: out <= 16'hFCD9;    16'd54057: out <= 16'hFDD9;    16'd54058: out <= 16'hFF27;    16'd54059: out <= 16'hFBD6;
    16'd54060: out <= 16'hFBE1;    16'd54061: out <= 16'hFBB0;    16'd54062: out <= 16'h0044;    16'd54063: out <= 16'h037F;
    16'd54064: out <= 16'h0964;    16'd54065: out <= 16'h03B5;    16'd54066: out <= 16'hFD85;    16'd54067: out <= 16'h0175;
    16'd54068: out <= 16'hFA87;    16'd54069: out <= 16'h0470;    16'd54070: out <= 16'h0D72;    16'd54071: out <= 16'h08C0;
    16'd54072: out <= 16'hFF6D;    16'd54073: out <= 16'h0DB3;    16'd54074: out <= 16'hF87A;    16'd54075: out <= 16'h01A8;
    16'd54076: out <= 16'h02F0;    16'd54077: out <= 16'hFDAA;    16'd54078: out <= 16'h0116;    16'd54079: out <= 16'h06AE;
    16'd54080: out <= 16'h0457;    16'd54081: out <= 16'h0569;    16'd54082: out <= 16'h02D1;    16'd54083: out <= 16'h0EDA;
    16'd54084: out <= 16'hFD70;    16'd54085: out <= 16'h073E;    16'd54086: out <= 16'h04A9;    16'd54087: out <= 16'h017C;
    16'd54088: out <= 16'h04D6;    16'd54089: out <= 16'h039F;    16'd54090: out <= 16'h0A01;    16'd54091: out <= 16'h0180;
    16'd54092: out <= 16'h0391;    16'd54093: out <= 16'h008B;    16'd54094: out <= 16'hFFC8;    16'd54095: out <= 16'h0C80;
    16'd54096: out <= 16'h083A;    16'd54097: out <= 16'h0592;    16'd54098: out <= 16'h02E3;    16'd54099: out <= 16'h051F;
    16'd54100: out <= 16'h0642;    16'd54101: out <= 16'hFB4A;    16'd54102: out <= 16'h0432;    16'd54103: out <= 16'h01C1;
    16'd54104: out <= 16'h0196;    16'd54105: out <= 16'h0268;    16'd54106: out <= 16'h06A2;    16'd54107: out <= 16'hFFC5;
    16'd54108: out <= 16'h0039;    16'd54109: out <= 16'h0712;    16'd54110: out <= 16'h0A3D;    16'd54111: out <= 16'hFECE;
    16'd54112: out <= 16'h0620;    16'd54113: out <= 16'hFCD3;    16'd54114: out <= 16'hFC69;    16'd54115: out <= 16'h02E1;
    16'd54116: out <= 16'hFF97;    16'd54117: out <= 16'hF853;    16'd54118: out <= 16'h0285;    16'd54119: out <= 16'hF6BF;
    16'd54120: out <= 16'hFC8E;    16'd54121: out <= 16'h06C8;    16'd54122: out <= 16'h0735;    16'd54123: out <= 16'hF5C0;
    16'd54124: out <= 16'hFE8F;    16'd54125: out <= 16'h03C7;    16'd54126: out <= 16'h0598;    16'd54127: out <= 16'hFFCC;
    16'd54128: out <= 16'hF6F9;    16'd54129: out <= 16'h06D3;    16'd54130: out <= 16'h014F;    16'd54131: out <= 16'h0091;
    16'd54132: out <= 16'h01E0;    16'd54133: out <= 16'hFFFF;    16'd54134: out <= 16'hFFD5;    16'd54135: out <= 16'hFDF5;
    16'd54136: out <= 16'hFEE0;    16'd54137: out <= 16'h03CF;    16'd54138: out <= 16'h064F;    16'd54139: out <= 16'hFD34;
    16'd54140: out <= 16'h0118;    16'd54141: out <= 16'h0BA8;    16'd54142: out <= 16'h02DE;    16'd54143: out <= 16'h0881;
    16'd54144: out <= 16'h0294;    16'd54145: out <= 16'h00C8;    16'd54146: out <= 16'h0442;    16'd54147: out <= 16'h00A0;
    16'd54148: out <= 16'h05B6;    16'd54149: out <= 16'h024B;    16'd54150: out <= 16'h092F;    16'd54151: out <= 16'h08B6;
    16'd54152: out <= 16'h098D;    16'd54153: out <= 16'h0409;    16'd54154: out <= 16'h041E;    16'd54155: out <= 16'h016A;
    16'd54156: out <= 16'h0349;    16'd54157: out <= 16'h0033;    16'd54158: out <= 16'h05A0;    16'd54159: out <= 16'h0864;
    16'd54160: out <= 16'hFFAA;    16'd54161: out <= 16'h0571;    16'd54162: out <= 16'h031F;    16'd54163: out <= 16'h03A6;
    16'd54164: out <= 16'h0B94;    16'd54165: out <= 16'h03AF;    16'd54166: out <= 16'h005E;    16'd54167: out <= 16'h07A4;
    16'd54168: out <= 16'h04DE;    16'd54169: out <= 16'h073E;    16'd54170: out <= 16'h0667;    16'd54171: out <= 16'h0399;
    16'd54172: out <= 16'h04B9;    16'd54173: out <= 16'h050D;    16'd54174: out <= 16'h0892;    16'd54175: out <= 16'h08A7;
    16'd54176: out <= 16'h0279;    16'd54177: out <= 16'h0647;    16'd54178: out <= 16'h043B;    16'd54179: out <= 16'h07CC;
    16'd54180: out <= 16'h040D;    16'd54181: out <= 16'h07F6;    16'd54182: out <= 16'h0081;    16'd54183: out <= 16'h09A4;
    16'd54184: out <= 16'h0622;    16'd54185: out <= 16'h04C2;    16'd54186: out <= 16'h02A9;    16'd54187: out <= 16'h01A8;
    16'd54188: out <= 16'h09F4;    16'd54189: out <= 16'h0338;    16'd54190: out <= 16'h0B39;    16'd54191: out <= 16'h0651;
    16'd54192: out <= 16'h0311;    16'd54193: out <= 16'h0A3F;    16'd54194: out <= 16'h0859;    16'd54195: out <= 16'hFC91;
    16'd54196: out <= 16'h08F3;    16'd54197: out <= 16'hFE30;    16'd54198: out <= 16'h046D;    16'd54199: out <= 16'h012C;
    16'd54200: out <= 16'h0546;    16'd54201: out <= 16'h0B1C;    16'd54202: out <= 16'h09DC;    16'd54203: out <= 16'h08B9;
    16'd54204: out <= 16'hFF6F;    16'd54205: out <= 16'h04AB;    16'd54206: out <= 16'h05FA;    16'd54207: out <= 16'h0834;
    16'd54208: out <= 16'h068E;    16'd54209: out <= 16'h0743;    16'd54210: out <= 16'h0453;    16'd54211: out <= 16'hF68E;
    16'd54212: out <= 16'h0549;    16'd54213: out <= 16'hFEB1;    16'd54214: out <= 16'hF8C5;    16'd54215: out <= 16'h0011;
    16'd54216: out <= 16'h0028;    16'd54217: out <= 16'h019E;    16'd54218: out <= 16'hFB5A;    16'd54219: out <= 16'h0493;
    16'd54220: out <= 16'hFBD7;    16'd54221: out <= 16'h0184;    16'd54222: out <= 16'hFE16;    16'd54223: out <= 16'hFE4E;
    16'd54224: out <= 16'h06B1;    16'd54225: out <= 16'h0686;    16'd54226: out <= 16'h02C5;    16'd54227: out <= 16'h0142;
    16'd54228: out <= 16'hFBA6;    16'd54229: out <= 16'hFDFF;    16'd54230: out <= 16'hFC3D;    16'd54231: out <= 16'hFE90;
    16'd54232: out <= 16'hFDE0;    16'd54233: out <= 16'h026E;    16'd54234: out <= 16'h0046;    16'd54235: out <= 16'hFF61;
    16'd54236: out <= 16'h028E;    16'd54237: out <= 16'h05DC;    16'd54238: out <= 16'h0568;    16'd54239: out <= 16'h0474;
    16'd54240: out <= 16'h07AF;    16'd54241: out <= 16'h03FD;    16'd54242: out <= 16'h00E3;    16'd54243: out <= 16'h044D;
    16'd54244: out <= 16'h00E8;    16'd54245: out <= 16'hFD1F;    16'd54246: out <= 16'h04A3;    16'd54247: out <= 16'h03AD;
    16'd54248: out <= 16'hF989;    16'd54249: out <= 16'h024E;    16'd54250: out <= 16'hFF8C;    16'd54251: out <= 16'hF8A1;
    16'd54252: out <= 16'hF870;    16'd54253: out <= 16'h0634;    16'd54254: out <= 16'hFFE5;    16'd54255: out <= 16'h04B0;
    16'd54256: out <= 16'hFD94;    16'd54257: out <= 16'hFEF7;    16'd54258: out <= 16'hFB8C;    16'd54259: out <= 16'hFB96;
    16'd54260: out <= 16'h004C;    16'd54261: out <= 16'hFD25;    16'd54262: out <= 16'hFF6F;    16'd54263: out <= 16'h04AB;
    16'd54264: out <= 16'h02CD;    16'd54265: out <= 16'h018B;    16'd54266: out <= 16'h02D8;    16'd54267: out <= 16'hFDB9;
    16'd54268: out <= 16'hFDB2;    16'd54269: out <= 16'h03A6;    16'd54270: out <= 16'hFFF1;    16'd54271: out <= 16'hFB83;
    16'd54272: out <= 16'h0372;    16'd54273: out <= 16'hFFFD;    16'd54274: out <= 16'h0261;    16'd54275: out <= 16'hFFCD;
    16'd54276: out <= 16'h01C7;    16'd54277: out <= 16'h0080;    16'd54278: out <= 16'hFE3C;    16'd54279: out <= 16'hFF9E;
    16'd54280: out <= 16'hFB1A;    16'd54281: out <= 16'hFEBF;    16'd54282: out <= 16'h0250;    16'd54283: out <= 16'hFF90;
    16'd54284: out <= 16'h01CB;    16'd54285: out <= 16'hFD18;    16'd54286: out <= 16'hFF97;    16'd54287: out <= 16'hF814;
    16'd54288: out <= 16'h00E1;    16'd54289: out <= 16'hFD7D;    16'd54290: out <= 16'h02B1;    16'd54291: out <= 16'h037E;
    16'd54292: out <= 16'h0130;    16'd54293: out <= 16'hFF1F;    16'd54294: out <= 16'h019A;    16'd54295: out <= 16'hFA2C;
    16'd54296: out <= 16'hF9C7;    16'd54297: out <= 16'hF6CC;    16'd54298: out <= 16'hFF80;    16'd54299: out <= 16'hFFB1;
    16'd54300: out <= 16'hF98A;    16'd54301: out <= 16'hFED9;    16'd54302: out <= 16'hFD38;    16'd54303: out <= 16'h01B2;
    16'd54304: out <= 16'h002F;    16'd54305: out <= 16'hFA7F;    16'd54306: out <= 16'h0235;    16'd54307: out <= 16'hFF3F;
    16'd54308: out <= 16'hFCBC;    16'd54309: out <= 16'hFF50;    16'd54310: out <= 16'hFED3;    16'd54311: out <= 16'h0251;
    16'd54312: out <= 16'h006F;    16'd54313: out <= 16'h0113;    16'd54314: out <= 16'h0454;    16'd54315: out <= 16'h06F4;
    16'd54316: out <= 16'h0552;    16'd54317: out <= 16'h0296;    16'd54318: out <= 16'h0146;    16'd54319: out <= 16'hFA35;
    16'd54320: out <= 16'h056F;    16'd54321: out <= 16'hFF52;    16'd54322: out <= 16'h00F8;    16'd54323: out <= 16'h02A8;
    16'd54324: out <= 16'h0502;    16'd54325: out <= 16'h0219;    16'd54326: out <= 16'hFF30;    16'd54327: out <= 16'h0648;
    16'd54328: out <= 16'h0691;    16'd54329: out <= 16'hFFE3;    16'd54330: out <= 16'h04B5;    16'd54331: out <= 16'h05B9;
    16'd54332: out <= 16'h02A8;    16'd54333: out <= 16'h04D8;    16'd54334: out <= 16'h078B;    16'd54335: out <= 16'h0A48;
    16'd54336: out <= 16'h0546;    16'd54337: out <= 16'h06A2;    16'd54338: out <= 16'h05CD;    16'd54339: out <= 16'hFF0C;
    16'd54340: out <= 16'h00B1;    16'd54341: out <= 16'h065D;    16'd54342: out <= 16'h02DA;    16'd54343: out <= 16'h0822;
    16'd54344: out <= 16'h07A2;    16'd54345: out <= 16'h032A;    16'd54346: out <= 16'h06B9;    16'd54347: out <= 16'h021E;
    16'd54348: out <= 16'hFF9A;    16'd54349: out <= 16'h058F;    16'd54350: out <= 16'h01A4;    16'd54351: out <= 16'hFC0D;
    16'd54352: out <= 16'hFED9;    16'd54353: out <= 16'h026B;    16'd54354: out <= 16'h047C;    16'd54355: out <= 16'h039B;
    16'd54356: out <= 16'h0C62;    16'd54357: out <= 16'hFF9D;    16'd54358: out <= 16'hFFEC;    16'd54359: out <= 16'h03C5;
    16'd54360: out <= 16'h0820;    16'd54361: out <= 16'h01E1;    16'd54362: out <= 16'h071F;    16'd54363: out <= 16'h029B;
    16'd54364: out <= 16'h03B0;    16'd54365: out <= 16'h0651;    16'd54366: out <= 16'h01C6;    16'd54367: out <= 16'h069D;
    16'd54368: out <= 16'hFEA4;    16'd54369: out <= 16'hFD89;    16'd54370: out <= 16'hFF29;    16'd54371: out <= 16'hFDE7;
    16'd54372: out <= 16'h043D;    16'd54373: out <= 16'hFEF7;    16'd54374: out <= 16'hFE40;    16'd54375: out <= 16'hFF9C;
    16'd54376: out <= 16'h0211;    16'd54377: out <= 16'hFB2C;    16'd54378: out <= 16'h03E2;    16'd54379: out <= 16'hFDD7;
    16'd54380: out <= 16'hFFD3;    16'd54381: out <= 16'h03D0;    16'd54382: out <= 16'hFBA3;    16'd54383: out <= 16'h0183;
    16'd54384: out <= 16'h0275;    16'd54385: out <= 16'h03D7;    16'd54386: out <= 16'hFF70;    16'd54387: out <= 16'h0486;
    16'd54388: out <= 16'h01B8;    16'd54389: out <= 16'h011E;    16'd54390: out <= 16'hFEEC;    16'd54391: out <= 16'hFF5A;
    16'd54392: out <= 16'h012E;    16'd54393: out <= 16'h0319;    16'd54394: out <= 16'hFCDE;    16'd54395: out <= 16'hFC90;
    16'd54396: out <= 16'hFF4B;    16'd54397: out <= 16'h0345;    16'd54398: out <= 16'h00E8;    16'd54399: out <= 16'hFAF7;
    16'd54400: out <= 16'h026C;    16'd54401: out <= 16'hFE36;    16'd54402: out <= 16'hFEB1;    16'd54403: out <= 16'h040A;
    16'd54404: out <= 16'h06DE;    16'd54405: out <= 16'h052D;    16'd54406: out <= 16'hFECD;    16'd54407: out <= 16'h02BF;
    16'd54408: out <= 16'hFD6D;    16'd54409: out <= 16'h0128;    16'd54410: out <= 16'hFFC4;    16'd54411: out <= 16'h0567;
    16'd54412: out <= 16'h04FC;    16'd54413: out <= 16'h01F1;    16'd54414: out <= 16'h04AA;    16'd54415: out <= 16'h07EE;
    16'd54416: out <= 16'hFFD5;    16'd54417: out <= 16'h01D0;    16'd54418: out <= 16'h066E;    16'd54419: out <= 16'h0450;
    16'd54420: out <= 16'h0634;    16'd54421: out <= 16'h01FF;    16'd54422: out <= 16'h0581;    16'd54423: out <= 16'h095D;
    16'd54424: out <= 16'h064D;    16'd54425: out <= 16'hFAE9;    16'd54426: out <= 16'h044B;    16'd54427: out <= 16'h0074;
    16'd54428: out <= 16'h02A1;    16'd54429: out <= 16'h0074;    16'd54430: out <= 16'h02C8;    16'd54431: out <= 16'hFAEF;
    16'd54432: out <= 16'h0558;    16'd54433: out <= 16'h03AC;    16'd54434: out <= 16'h06BB;    16'd54435: out <= 16'hFD24;
    16'd54436: out <= 16'h0214;    16'd54437: out <= 16'h0638;    16'd54438: out <= 16'h09E0;    16'd54439: out <= 16'h062E;
    16'd54440: out <= 16'h08E9;    16'd54441: out <= 16'h085A;    16'd54442: out <= 16'h02BD;    16'd54443: out <= 16'h035C;
    16'd54444: out <= 16'h05CB;    16'd54445: out <= 16'h0243;    16'd54446: out <= 16'h032F;    16'd54447: out <= 16'h021B;
    16'd54448: out <= 16'h0789;    16'd54449: out <= 16'h0405;    16'd54450: out <= 16'h0351;    16'd54451: out <= 16'h01C5;
    16'd54452: out <= 16'h02D4;    16'd54453: out <= 16'h01FB;    16'd54454: out <= 16'h0896;    16'd54455: out <= 16'h06B0;
    16'd54456: out <= 16'h0747;    16'd54457: out <= 16'h0213;    16'd54458: out <= 16'h0588;    16'd54459: out <= 16'h06AA;
    16'd54460: out <= 16'h058D;    16'd54461: out <= 16'h08D4;    16'd54462: out <= 16'h0219;    16'd54463: out <= 16'h00E9;
    16'd54464: out <= 16'h0331;    16'd54465: out <= 16'h0426;    16'd54466: out <= 16'h0548;    16'd54467: out <= 16'hFEE8;
    16'd54468: out <= 16'h0001;    16'd54469: out <= 16'h01F4;    16'd54470: out <= 16'hF984;    16'd54471: out <= 16'hFB61;
    16'd54472: out <= 16'h0647;    16'd54473: out <= 16'hFA73;    16'd54474: out <= 16'h058F;    16'd54475: out <= 16'hFF95;
    16'd54476: out <= 16'h03B7;    16'd54477: out <= 16'h018C;    16'd54478: out <= 16'h03A7;    16'd54479: out <= 16'hF73B;
    16'd54480: out <= 16'hFC0B;    16'd54481: out <= 16'hFC15;    16'd54482: out <= 16'h08B9;    16'd54483: out <= 16'hFF40;
    16'd54484: out <= 16'h03A6;    16'd54485: out <= 16'hFF80;    16'd54486: out <= 16'h0317;    16'd54487: out <= 16'h0596;
    16'd54488: out <= 16'hF932;    16'd54489: out <= 16'h001F;    16'd54490: out <= 16'h06B4;    16'd54491: out <= 16'hFC25;
    16'd54492: out <= 16'h0233;    16'd54493: out <= 16'hFF9C;    16'd54494: out <= 16'h06A9;    16'd54495: out <= 16'h0585;
    16'd54496: out <= 16'h00E4;    16'd54497: out <= 16'h0169;    16'd54498: out <= 16'hF7C1;    16'd54499: out <= 16'h0379;
    16'd54500: out <= 16'hF970;    16'd54501: out <= 16'hFF44;    16'd54502: out <= 16'h0026;    16'd54503: out <= 16'hFC80;
    16'd54504: out <= 16'hFB85;    16'd54505: out <= 16'hFF27;    16'd54506: out <= 16'h0773;    16'd54507: out <= 16'hFF19;
    16'd54508: out <= 16'h03E0;    16'd54509: out <= 16'hFCC3;    16'd54510: out <= 16'h04B7;    16'd54511: out <= 16'h0197;
    16'd54512: out <= 16'h03CA;    16'd54513: out <= 16'hFD51;    16'd54514: out <= 16'h0193;    16'd54515: out <= 16'hFD61;
    16'd54516: out <= 16'h0010;    16'd54517: out <= 16'hFDB3;    16'd54518: out <= 16'hFA4A;    16'd54519: out <= 16'h064D;
    16'd54520: out <= 16'hFDDE;    16'd54521: out <= 16'h05C5;    16'd54522: out <= 16'h02EF;    16'd54523: out <= 16'h0200;
    16'd54524: out <= 16'h0089;    16'd54525: out <= 16'h000D;    16'd54526: out <= 16'hFCEA;    16'd54527: out <= 16'h06C2;
    16'd54528: out <= 16'h02DE;    16'd54529: out <= 16'hFF16;    16'd54530: out <= 16'h0221;    16'd54531: out <= 16'hFF30;
    16'd54532: out <= 16'h0054;    16'd54533: out <= 16'hFF07;    16'd54534: out <= 16'h0840;    16'd54535: out <= 16'h043C;
    16'd54536: out <= 16'hFBB4;    16'd54537: out <= 16'hFFCA;    16'd54538: out <= 16'hFF29;    16'd54539: out <= 16'hFBB0;
    16'd54540: out <= 16'hFD4B;    16'd54541: out <= 16'h010B;    16'd54542: out <= 16'hF9FB;    16'd54543: out <= 16'hFEFB;
    16'd54544: out <= 16'h053D;    16'd54545: out <= 16'h029A;    16'd54546: out <= 16'h0005;    16'd54547: out <= 16'h0498;
    16'd54548: out <= 16'h0213;    16'd54549: out <= 16'hF8BB;    16'd54550: out <= 16'h00AE;    16'd54551: out <= 16'h0433;
    16'd54552: out <= 16'hFB78;    16'd54553: out <= 16'hFB15;    16'd54554: out <= 16'h07D6;    16'd54555: out <= 16'h0497;
    16'd54556: out <= 16'hFBDF;    16'd54557: out <= 16'hF7DE;    16'd54558: out <= 16'hFA56;    16'd54559: out <= 16'hF9A6;
    16'd54560: out <= 16'h00B6;    16'd54561: out <= 16'h0037;    16'd54562: out <= 16'hFCA4;    16'd54563: out <= 16'h011B;
    16'd54564: out <= 16'hFB84;    16'd54565: out <= 16'h0107;    16'd54566: out <= 16'h02B1;    16'd54567: out <= 16'hFE1B;
    16'd54568: out <= 16'h0038;    16'd54569: out <= 16'hFDF5;    16'd54570: out <= 16'hFBCA;    16'd54571: out <= 16'hFD1E;
    16'd54572: out <= 16'h05F5;    16'd54573: out <= 16'hFAF9;    16'd54574: out <= 16'hFEBE;    16'd54575: out <= 16'hFED1;
    16'd54576: out <= 16'h03A7;    16'd54577: out <= 16'h05AD;    16'd54578: out <= 16'h062F;    16'd54579: out <= 16'hFE77;
    16'd54580: out <= 16'hFDA3;    16'd54581: out <= 16'h00E0;    16'd54582: out <= 16'h0373;    16'd54583: out <= 16'h05B7;
    16'd54584: out <= 16'h03D5;    16'd54585: out <= 16'h067F;    16'd54586: out <= 16'h084F;    16'd54587: out <= 16'h0190;
    16'd54588: out <= 16'h00B7;    16'd54589: out <= 16'hFED8;    16'd54590: out <= 16'h0620;    16'd54591: out <= 16'hFAD8;
    16'd54592: out <= 16'h03CE;    16'd54593: out <= 16'h0926;    16'd54594: out <= 16'h0671;    16'd54595: out <= 16'h03F7;
    16'd54596: out <= 16'hFAF1;    16'd54597: out <= 16'h02C7;    16'd54598: out <= 16'hFEF7;    16'd54599: out <= 16'h03D6;
    16'd54600: out <= 16'h017B;    16'd54601: out <= 16'h071C;    16'd54602: out <= 16'h0955;    16'd54603: out <= 16'h056B;
    16'd54604: out <= 16'h0285;    16'd54605: out <= 16'h061B;    16'd54606: out <= 16'h0560;    16'd54607: out <= 16'h03E1;
    16'd54608: out <= 16'h061A;    16'd54609: out <= 16'h0555;    16'd54610: out <= 16'h078F;    16'd54611: out <= 16'h02CD;
    16'd54612: out <= 16'h0739;    16'd54613: out <= 16'h0370;    16'd54614: out <= 16'h018B;    16'd54615: out <= 16'h05ED;
    16'd54616: out <= 16'hF9C2;    16'd54617: out <= 16'h0165;    16'd54618: out <= 16'h05C6;    16'd54619: out <= 16'h04B8;
    16'd54620: out <= 16'hFEE4;    16'd54621: out <= 16'h031E;    16'd54622: out <= 16'h07C7;    16'd54623: out <= 16'h0778;
    16'd54624: out <= 16'h0098;    16'd54625: out <= 16'h0A21;    16'd54626: out <= 16'hFF2A;    16'd54627: out <= 16'h03F0;
    16'd54628: out <= 16'h084B;    16'd54629: out <= 16'h020D;    16'd54630: out <= 16'hFAD2;    16'd54631: out <= 16'hFE41;
    16'd54632: out <= 16'h0012;    16'd54633: out <= 16'h0228;    16'd54634: out <= 16'hF914;    16'd54635: out <= 16'h01D8;
    16'd54636: out <= 16'hFEF2;    16'd54637: out <= 16'h02AF;    16'd54638: out <= 16'h042E;    16'd54639: out <= 16'h0568;
    16'd54640: out <= 16'h046B;    16'd54641: out <= 16'h0A2A;    16'd54642: out <= 16'h073D;    16'd54643: out <= 16'h051E;
    16'd54644: out <= 16'h0610;    16'd54645: out <= 16'hFCD9;    16'd54646: out <= 16'h0332;    16'd54647: out <= 16'h05BD;
    16'd54648: out <= 16'h0533;    16'd54649: out <= 16'hFE46;    16'd54650: out <= 16'h0363;    16'd54651: out <= 16'h07C5;
    16'd54652: out <= 16'h06D2;    16'd54653: out <= 16'h0412;    16'd54654: out <= 16'h0771;    16'd54655: out <= 16'h057A;
    16'd54656: out <= 16'h03E4;    16'd54657: out <= 16'h05CF;    16'd54658: out <= 16'h01AE;    16'd54659: out <= 16'h07E1;
    16'd54660: out <= 16'h0594;    16'd54661: out <= 16'hFF06;    16'd54662: out <= 16'h0401;    16'd54663: out <= 16'h02A9;
    16'd54664: out <= 16'h0431;    16'd54665: out <= 16'h0574;    16'd54666: out <= 16'h057A;    16'd54667: out <= 16'h0482;
    16'd54668: out <= 16'hFFA1;    16'd54669: out <= 16'h0A4C;    16'd54670: out <= 16'h065F;    16'd54671: out <= 16'h015B;
    16'd54672: out <= 16'h0C39;    16'd54673: out <= 16'h005C;    16'd54674: out <= 16'h04A9;    16'd54675: out <= 16'hFF2D;
    16'd54676: out <= 16'h028C;    16'd54677: out <= 16'h01A0;    16'd54678: out <= 16'hF9D4;    16'd54679: out <= 16'h080E;
    16'd54680: out <= 16'hFFA5;    16'd54681: out <= 16'h0B2F;    16'd54682: out <= 16'h057A;    16'd54683: out <= 16'h0726;
    16'd54684: out <= 16'h03A0;    16'd54685: out <= 16'hFE39;    16'd54686: out <= 16'hFC0C;    16'd54687: out <= 16'hFB3E;
    16'd54688: out <= 16'h02CA;    16'd54689: out <= 16'h05A8;    16'd54690: out <= 16'h05BC;    16'd54691: out <= 16'h048B;
    16'd54692: out <= 16'h0449;    16'd54693: out <= 16'hFF92;    16'd54694: out <= 16'h0849;    16'd54695: out <= 16'hFB7D;
    16'd54696: out <= 16'h0275;    16'd54697: out <= 16'h0824;    16'd54698: out <= 16'h04F4;    16'd54699: out <= 16'h0842;
    16'd54700: out <= 16'h0573;    16'd54701: out <= 16'hF959;    16'd54702: out <= 16'h0077;    16'd54703: out <= 16'hFED5;
    16'd54704: out <= 16'h1072;    16'd54705: out <= 16'h0315;    16'd54706: out <= 16'h06FE;    16'd54707: out <= 16'h04FE;
    16'd54708: out <= 16'h05C5;    16'd54709: out <= 16'h05FD;    16'd54710: out <= 16'h0585;    16'd54711: out <= 16'hFFB3;
    16'd54712: out <= 16'h059D;    16'd54713: out <= 16'h0304;    16'd54714: out <= 16'h014C;    16'd54715: out <= 16'hFFEF;
    16'd54716: out <= 16'h01DB;    16'd54717: out <= 16'h00EE;    16'd54718: out <= 16'h0431;    16'd54719: out <= 16'hF9E5;
    16'd54720: out <= 16'h02F2;    16'd54721: out <= 16'h07D5;    16'd54722: out <= 16'hFF0E;    16'd54723: out <= 16'h05BD;
    16'd54724: out <= 16'h02AD;    16'd54725: out <= 16'h0293;    16'd54726: out <= 16'h0859;    16'd54727: out <= 16'h01D2;
    16'd54728: out <= 16'hFCC9;    16'd54729: out <= 16'hFE92;    16'd54730: out <= 16'h041D;    16'd54731: out <= 16'hFDE3;
    16'd54732: out <= 16'h03B8;    16'd54733: out <= 16'h07A0;    16'd54734: out <= 16'h06C4;    16'd54735: out <= 16'hFFDB;
    16'd54736: out <= 16'h03CC;    16'd54737: out <= 16'h0007;    16'd54738: out <= 16'h00A7;    16'd54739: out <= 16'h0191;
    16'd54740: out <= 16'h014B;    16'd54741: out <= 16'hF8DF;    16'd54742: out <= 16'h0292;    16'd54743: out <= 16'hFAE1;
    16'd54744: out <= 16'hFE13;    16'd54745: out <= 16'h04EF;    16'd54746: out <= 16'hFE50;    16'd54747: out <= 16'h0460;
    16'd54748: out <= 16'h0401;    16'd54749: out <= 16'h003C;    16'd54750: out <= 16'hFFA2;    16'd54751: out <= 16'h0423;
    16'd54752: out <= 16'h083E;    16'd54753: out <= 16'hFE3A;    16'd54754: out <= 16'h0093;    16'd54755: out <= 16'h0259;
    16'd54756: out <= 16'h0595;    16'd54757: out <= 16'h021D;    16'd54758: out <= 16'hFC5E;    16'd54759: out <= 16'hFFD1;
    16'd54760: out <= 16'hFA7A;    16'd54761: out <= 16'hFB89;    16'd54762: out <= 16'hFFCA;    16'd54763: out <= 16'hFBAE;
    16'd54764: out <= 16'hFB71;    16'd54765: out <= 16'h02E6;    16'd54766: out <= 16'hF9D2;    16'd54767: out <= 16'hFDD5;
    16'd54768: out <= 16'hFFE2;    16'd54769: out <= 16'h00DC;    16'd54770: out <= 16'h0076;    16'd54771: out <= 16'h0150;
    16'd54772: out <= 16'h0326;    16'd54773: out <= 16'h0046;    16'd54774: out <= 16'h0839;    16'd54775: out <= 16'h056F;
    16'd54776: out <= 16'h0036;    16'd54777: out <= 16'h026D;    16'd54778: out <= 16'h03E8;    16'd54779: out <= 16'hFB54;
    16'd54780: out <= 16'h0DD2;    16'd54781: out <= 16'hFD02;    16'd54782: out <= 16'hF4E5;    16'd54783: out <= 16'hFA20;
    16'd54784: out <= 16'hFC9E;    16'd54785: out <= 16'hFE7D;    16'd54786: out <= 16'h0202;    16'd54787: out <= 16'h0678;
    16'd54788: out <= 16'hFDC4;    16'd54789: out <= 16'hF8AC;    16'd54790: out <= 16'hFAE2;    16'd54791: out <= 16'h05C7;
    16'd54792: out <= 16'h016A;    16'd54793: out <= 16'h009C;    16'd54794: out <= 16'h04ED;    16'd54795: out <= 16'h0371;
    16'd54796: out <= 16'h02B5;    16'd54797: out <= 16'hFE8C;    16'd54798: out <= 16'h02D8;    16'd54799: out <= 16'hF9F4;
    16'd54800: out <= 16'h02EF;    16'd54801: out <= 16'h0100;    16'd54802: out <= 16'h04E6;    16'd54803: out <= 16'h011F;
    16'd54804: out <= 16'hFE74;    16'd54805: out <= 16'h027A;    16'd54806: out <= 16'hFADA;    16'd54807: out <= 16'h0163;
    16'd54808: out <= 16'hFD41;    16'd54809: out <= 16'h0194;    16'd54810: out <= 16'hFF3C;    16'd54811: out <= 16'hFEDF;
    16'd54812: out <= 16'hFFB2;    16'd54813: out <= 16'hFD7C;    16'd54814: out <= 16'hF9B3;    16'd54815: out <= 16'hFD98;
    16'd54816: out <= 16'hF940;    16'd54817: out <= 16'hFEEA;    16'd54818: out <= 16'h077E;    16'd54819: out <= 16'hFE5B;
    16'd54820: out <= 16'h0396;    16'd54821: out <= 16'h0441;    16'd54822: out <= 16'hFBD4;    16'd54823: out <= 16'hFA4B;
    16'd54824: out <= 16'hFD43;    16'd54825: out <= 16'h04F3;    16'd54826: out <= 16'hFFF2;    16'd54827: out <= 16'h0481;
    16'd54828: out <= 16'h0129;    16'd54829: out <= 16'h00F8;    16'd54830: out <= 16'h01FF;    16'd54831: out <= 16'hFDB5;
    16'd54832: out <= 16'h00AB;    16'd54833: out <= 16'hFDCD;    16'd54834: out <= 16'h03FE;    16'd54835: out <= 16'h0221;
    16'd54836: out <= 16'hFEF9;    16'd54837: out <= 16'hFF05;    16'd54838: out <= 16'h069E;    16'd54839: out <= 16'h0C38;
    16'd54840: out <= 16'h06B3;    16'd54841: out <= 16'h0834;    16'd54842: out <= 16'h061E;    16'd54843: out <= 16'hFFEC;
    16'd54844: out <= 16'h051D;    16'd54845: out <= 16'h02EB;    16'd54846: out <= 16'h0185;    16'd54847: out <= 16'h077F;
    16'd54848: out <= 16'h00F1;    16'd54849: out <= 16'h0A03;    16'd54850: out <= 16'h05EF;    16'd54851: out <= 16'hFC36;
    16'd54852: out <= 16'h01E8;    16'd54853: out <= 16'h05A9;    16'd54854: out <= 16'h024B;    16'd54855: out <= 16'hFE56;
    16'd54856: out <= 16'h0A64;    16'd54857: out <= 16'h03D8;    16'd54858: out <= 16'h0341;    16'd54859: out <= 16'h0057;
    16'd54860: out <= 16'h0500;    16'd54861: out <= 16'h04D4;    16'd54862: out <= 16'h0184;    16'd54863: out <= 16'h0162;
    16'd54864: out <= 16'h08AA;    16'd54865: out <= 16'h09F1;    16'd54866: out <= 16'h0961;    16'd54867: out <= 16'h002F;
    16'd54868: out <= 16'h01C8;    16'd54869: out <= 16'h00FD;    16'd54870: out <= 16'h042F;    16'd54871: out <= 16'hFE07;
    16'd54872: out <= 16'h00DC;    16'd54873: out <= 16'h041F;    16'd54874: out <= 16'hFD85;    16'd54875: out <= 16'h03A1;
    16'd54876: out <= 16'h07A8;    16'd54877: out <= 16'h010D;    16'd54878: out <= 16'h0024;    16'd54879: out <= 16'h042C;
    16'd54880: out <= 16'h076E;    16'd54881: out <= 16'h02D9;    16'd54882: out <= 16'h0BC3;    16'd54883: out <= 16'h05E8;
    16'd54884: out <= 16'hFE9F;    16'd54885: out <= 16'h0A0B;    16'd54886: out <= 16'h02E5;    16'd54887: out <= 16'h01CE;
    16'd54888: out <= 16'h0174;    16'd54889: out <= 16'hFE8C;    16'd54890: out <= 16'h01E2;    16'd54891: out <= 16'h00DF;
    16'd54892: out <= 16'h02B3;    16'd54893: out <= 16'hFE8D;    16'd54894: out <= 16'h0498;    16'd54895: out <= 16'h00D0;
    16'd54896: out <= 16'h0755;    16'd54897: out <= 16'h03BC;    16'd54898: out <= 16'h07E6;    16'd54899: out <= 16'h04CA;
    16'd54900: out <= 16'h0A8E;    16'd54901: out <= 16'h0130;    16'd54902: out <= 16'h0530;    16'd54903: out <= 16'h0695;
    16'd54904: out <= 16'h0B3F;    16'd54905: out <= 16'h02A2;    16'd54906: out <= 16'h0468;    16'd54907: out <= 16'h0718;
    16'd54908: out <= 16'h01C7;    16'd54909: out <= 16'h02EA;    16'd54910: out <= 16'hFDF1;    16'd54911: out <= 16'h081D;
    16'd54912: out <= 16'h065B;    16'd54913: out <= 16'h0021;    16'd54914: out <= 16'h02F1;    16'd54915: out <= 16'h0693;
    16'd54916: out <= 16'h07C1;    16'd54917: out <= 16'h0358;    16'd54918: out <= 16'h0472;    16'd54919: out <= 16'h0818;
    16'd54920: out <= 16'h04F6;    16'd54921: out <= 16'h1097;    16'd54922: out <= 16'h11D2;    16'd54923: out <= 16'h006F;
    16'd54924: out <= 16'h02E3;    16'd54925: out <= 16'hFE29;    16'd54926: out <= 16'h08C0;    16'd54927: out <= 16'h0840;
    16'd54928: out <= 16'h0101;    16'd54929: out <= 16'h0251;    16'd54930: out <= 16'hFE78;    16'd54931: out <= 16'hFF41;
    16'd54932: out <= 16'hFDC8;    16'd54933: out <= 16'h0BBF;    16'd54934: out <= 16'hFDE4;    16'd54935: out <= 16'h0513;
    16'd54936: out <= 16'h0162;    16'd54937: out <= 16'hFE88;    16'd54938: out <= 16'h069A;    16'd54939: out <= 16'h00AA;
    16'd54940: out <= 16'h0D46;    16'd54941: out <= 16'h093C;    16'd54942: out <= 16'h07E6;    16'd54943: out <= 16'h0A98;
    16'd54944: out <= 16'h01BC;    16'd54945: out <= 16'h0555;    16'd54946: out <= 16'h03EF;    16'd54947: out <= 16'h057E;
    16'd54948: out <= 16'h00F1;    16'd54949: out <= 16'h0797;    16'd54950: out <= 16'h0552;    16'd54951: out <= 16'h0605;
    16'd54952: out <= 16'h0304;    16'd54953: out <= 16'h0450;    16'd54954: out <= 16'h06CF;    16'd54955: out <= 16'h07D4;
    16'd54956: out <= 16'hFB12;    16'd54957: out <= 16'h04C9;    16'd54958: out <= 16'h00F8;    16'd54959: out <= 16'h070D;
    16'd54960: out <= 16'hFF67;    16'd54961: out <= 16'hFE63;    16'd54962: out <= 16'h0946;    16'd54963: out <= 16'h03A9;
    16'd54964: out <= 16'h0623;    16'd54965: out <= 16'h021B;    16'd54966: out <= 16'h079A;    16'd54967: out <= 16'h03D7;
    16'd54968: out <= 16'h08C0;    16'd54969: out <= 16'h05D5;    16'd54970: out <= 16'h061F;    16'd54971: out <= 16'hFF8B;
    16'd54972: out <= 16'h05F9;    16'd54973: out <= 16'h02EE;    16'd54974: out <= 16'h0778;    16'd54975: out <= 16'h0598;
    16'd54976: out <= 16'h068C;    16'd54977: out <= 16'h012D;    16'd54978: out <= 16'h05E1;    16'd54979: out <= 16'h0172;
    16'd54980: out <= 16'hFD77;    16'd54981: out <= 16'hFF9A;    16'd54982: out <= 16'h01FD;    16'd54983: out <= 16'h01D4;
    16'd54984: out <= 16'hFAD6;    16'd54985: out <= 16'h0168;    16'd54986: out <= 16'hF8C2;    16'd54987: out <= 16'hFB1B;
    16'd54988: out <= 16'h0003;    16'd54989: out <= 16'h0286;    16'd54990: out <= 16'h061B;    16'd54991: out <= 16'h00D6;
    16'd54992: out <= 16'h02F0;    16'd54993: out <= 16'hFD25;    16'd54994: out <= 16'h0238;    16'd54995: out <= 16'h0132;
    16'd54996: out <= 16'hFF7A;    16'd54997: out <= 16'h0129;    16'd54998: out <= 16'h0015;    16'd54999: out <= 16'h050A;
    16'd55000: out <= 16'hFAFE;    16'd55001: out <= 16'hFCB0;    16'd55002: out <= 16'hFE26;    16'd55003: out <= 16'hF9DF;
    16'd55004: out <= 16'h0108;    16'd55005: out <= 16'h02B0;    16'd55006: out <= 16'h00C3;    16'd55007: out <= 16'h00DD;
    16'd55008: out <= 16'h014B;    16'd55009: out <= 16'h00CE;    16'd55010: out <= 16'hFF67;    16'd55011: out <= 16'h04A8;
    16'd55012: out <= 16'hFB76;    16'd55013: out <= 16'h0062;    16'd55014: out <= 16'hFAA8;    16'd55015: out <= 16'hFE07;
    16'd55016: out <= 16'h08C9;    16'd55017: out <= 16'hFD13;    16'd55018: out <= 16'h01A2;    16'd55019: out <= 16'hFA28;
    16'd55020: out <= 16'hFD5F;    16'd55021: out <= 16'hFD2B;    16'd55022: out <= 16'hFB6A;    16'd55023: out <= 16'h013D;
    16'd55024: out <= 16'h03C8;    16'd55025: out <= 16'h01AE;    16'd55026: out <= 16'hFBE6;    16'd55027: out <= 16'hFF61;
    16'd55028: out <= 16'h027F;    16'd55029: out <= 16'hFC6E;    16'd55030: out <= 16'hFCB4;    16'd55031: out <= 16'hFAB2;
    16'd55032: out <= 16'hFACD;    16'd55033: out <= 16'h00B2;    16'd55034: out <= 16'h02F2;    16'd55035: out <= 16'hFC35;
    16'd55036: out <= 16'h00DD;    16'd55037: out <= 16'hFE4D;    16'd55038: out <= 16'h05D4;    16'd55039: out <= 16'hFEF7;
    16'd55040: out <= 16'hFCFE;    16'd55041: out <= 16'h036B;    16'd55042: out <= 16'h0166;    16'd55043: out <= 16'hFBFE;
    16'd55044: out <= 16'h02B3;    16'd55045: out <= 16'hF9F9;    16'd55046: out <= 16'h03A3;    16'd55047: out <= 16'hF9F4;
    16'd55048: out <= 16'h044E;    16'd55049: out <= 16'hFD1C;    16'd55050: out <= 16'h05A0;    16'd55051: out <= 16'h0147;
    16'd55052: out <= 16'hFBF0;    16'd55053: out <= 16'hFBD8;    16'd55054: out <= 16'h01A5;    16'd55055: out <= 16'h0721;
    16'd55056: out <= 16'hFD5F;    16'd55057: out <= 16'h049C;    16'd55058: out <= 16'h05E8;    16'd55059: out <= 16'h0008;
    16'd55060: out <= 16'h0446;    16'd55061: out <= 16'h065B;    16'd55062: out <= 16'hFDF9;    16'd55063: out <= 16'hFAF6;
    16'd55064: out <= 16'hFF35;    16'd55065: out <= 16'hFCF6;    16'd55066: out <= 16'hFDAF;    16'd55067: out <= 16'h0069;
    16'd55068: out <= 16'hF9BD;    16'd55069: out <= 16'hFFEE;    16'd55070: out <= 16'hFD1C;    16'd55071: out <= 16'h0199;
    16'd55072: out <= 16'h032A;    16'd55073: out <= 16'h026D;    16'd55074: out <= 16'hFFD3;    16'd55075: out <= 16'h0280;
    16'd55076: out <= 16'h06EF;    16'd55077: out <= 16'h0381;    16'd55078: out <= 16'h02CE;    16'd55079: out <= 16'hFC26;
    16'd55080: out <= 16'hFD37;    16'd55081: out <= 16'hFEA2;    16'd55082: out <= 16'hFC20;    16'd55083: out <= 16'hFE19;
    16'd55084: out <= 16'h0580;    16'd55085: out <= 16'h0272;    16'd55086: out <= 16'h04A2;    16'd55087: out <= 16'hFE57;
    16'd55088: out <= 16'h00E3;    16'd55089: out <= 16'h05D0;    16'd55090: out <= 16'h0859;    16'd55091: out <= 16'h0882;
    16'd55092: out <= 16'hFEED;    16'd55093: out <= 16'h0C9D;    16'd55094: out <= 16'h01E3;    16'd55095: out <= 16'hFF5E;
    16'd55096: out <= 16'h055F;    16'd55097: out <= 16'h0619;    16'd55098: out <= 16'h0640;    16'd55099: out <= 16'hFA19;
    16'd55100: out <= 16'hFDB6;    16'd55101: out <= 16'h01FF;    16'd55102: out <= 16'h02B6;    16'd55103: out <= 16'h0392;
    16'd55104: out <= 16'h0810;    16'd55105: out <= 16'h0274;    16'd55106: out <= 16'h04C4;    16'd55107: out <= 16'h072D;
    16'd55108: out <= 16'hFF94;    16'd55109: out <= 16'h0652;    16'd55110: out <= 16'h0905;    16'd55111: out <= 16'h001A;
    16'd55112: out <= 16'h05C3;    16'd55113: out <= 16'h01D0;    16'd55114: out <= 16'h0661;    16'd55115: out <= 16'h0589;
    16'd55116: out <= 16'h089D;    16'd55117: out <= 16'h037F;    16'd55118: out <= 16'h0B70;    16'd55119: out <= 16'h0736;
    16'd55120: out <= 16'h02E1;    16'd55121: out <= 16'h0637;    16'd55122: out <= 16'h0215;    16'd55123: out <= 16'h0387;
    16'd55124: out <= 16'h0592;    16'd55125: out <= 16'h04CA;    16'd55126: out <= 16'h051C;    16'd55127: out <= 16'h05E2;
    16'd55128: out <= 16'h0872;    16'd55129: out <= 16'h008D;    16'd55130: out <= 16'h0A7D;    16'd55131: out <= 16'h0407;
    16'd55132: out <= 16'hFC2D;    16'd55133: out <= 16'h0523;    16'd55134: out <= 16'hFBED;    16'd55135: out <= 16'h02CA;
    16'd55136: out <= 16'hFE8A;    16'd55137: out <= 16'h01AB;    16'd55138: out <= 16'h009F;    16'd55139: out <= 16'h0219;
    16'd55140: out <= 16'hFFC8;    16'd55141: out <= 16'h0521;    16'd55142: out <= 16'hFE66;    16'd55143: out <= 16'hFDE4;
    16'd55144: out <= 16'h02BC;    16'd55145: out <= 16'hFFAB;    16'd55146: out <= 16'h0246;    16'd55147: out <= 16'h053C;
    16'd55148: out <= 16'h038D;    16'd55149: out <= 16'h05DC;    16'd55150: out <= 16'hFFED;    16'd55151: out <= 16'h06B7;
    16'd55152: out <= 16'h068C;    16'd55153: out <= 16'h085B;    16'd55154: out <= 16'hFCE0;    16'd55155: out <= 16'h03DC;
    16'd55156: out <= 16'h0035;    16'd55157: out <= 16'h02A4;    16'd55158: out <= 16'h0364;    16'd55159: out <= 16'h00DD;
    16'd55160: out <= 16'h0018;    16'd55161: out <= 16'h06C9;    16'd55162: out <= 16'h042C;    16'd55163: out <= 16'h0407;
    16'd55164: out <= 16'h0BD5;    16'd55165: out <= 16'h033F;    16'd55166: out <= 16'h039C;    16'd55167: out <= 16'h04AD;
    16'd55168: out <= 16'h0880;    16'd55169: out <= 16'h043A;    16'd55170: out <= 16'h0599;    16'd55171: out <= 16'h02AB;
    16'd55172: out <= 16'h029F;    16'd55173: out <= 16'hFFDD;    16'd55174: out <= 16'h0943;    16'd55175: out <= 16'h04F0;
    16'd55176: out <= 16'h01F6;    16'd55177: out <= 16'h0923;    16'd55178: out <= 16'h03F2;    16'd55179: out <= 16'h0342;
    16'd55180: out <= 16'h03C0;    16'd55181: out <= 16'h0632;    16'd55182: out <= 16'h013A;    16'd55183: out <= 16'hFF70;
    16'd55184: out <= 16'h0041;    16'd55185: out <= 16'h04A8;    16'd55186: out <= 16'h004C;    16'd55187: out <= 16'h04D1;
    16'd55188: out <= 16'h0384;    16'd55189: out <= 16'h00E6;    16'd55190: out <= 16'h07EA;    16'd55191: out <= 16'h0767;
    16'd55192: out <= 16'hFBF9;    16'd55193: out <= 16'h05EE;    16'd55194: out <= 16'h02A5;    16'd55195: out <= 16'hFB7F;
    16'd55196: out <= 16'h0426;    16'd55197: out <= 16'h0006;    16'd55198: out <= 16'h044B;    16'd55199: out <= 16'h0508;
    16'd55200: out <= 16'hFDAA;    16'd55201: out <= 16'h0B43;    16'd55202: out <= 16'hFEC3;    16'd55203: out <= 16'hFF9D;
    16'd55204: out <= 16'h00C4;    16'd55205: out <= 16'h012F;    16'd55206: out <= 16'h0698;    16'd55207: out <= 16'hFDAB;
    16'd55208: out <= 16'h03B1;    16'd55209: out <= 16'h04FE;    16'd55210: out <= 16'h0108;    16'd55211: out <= 16'h0039;
    16'd55212: out <= 16'h0435;    16'd55213: out <= 16'h0D18;    16'd55214: out <= 16'h0238;    16'd55215: out <= 16'hFF60;
    16'd55216: out <= 16'h0873;    16'd55217: out <= 16'h092D;    16'd55218: out <= 16'h0B3E;    16'd55219: out <= 16'h00C3;
    16'd55220: out <= 16'h04EF;    16'd55221: out <= 16'h0778;    16'd55222: out <= 16'h03CC;    16'd55223: out <= 16'h0299;
    16'd55224: out <= 16'h0785;    16'd55225: out <= 16'h00C5;    16'd55226: out <= 16'h0655;    16'd55227: out <= 16'h0410;
    16'd55228: out <= 16'h00CB;    16'd55229: out <= 16'h0486;    16'd55230: out <= 16'h0549;    16'd55231: out <= 16'h052A;
    16'd55232: out <= 16'hFE6C;    16'd55233: out <= 16'h02AD;    16'd55234: out <= 16'h0265;    16'd55235: out <= 16'hFBE8;
    16'd55236: out <= 16'h00B2;    16'd55237: out <= 16'hF5D0;    16'd55238: out <= 16'h0044;    16'd55239: out <= 16'hFFBA;
    16'd55240: out <= 16'hF5D9;    16'd55241: out <= 16'h0199;    16'd55242: out <= 16'hF9A0;    16'd55243: out <= 16'hFD49;
    16'd55244: out <= 16'h07CD;    16'd55245: out <= 16'hFD7C;    16'd55246: out <= 16'hFD18;    16'd55247: out <= 16'h01AC;
    16'd55248: out <= 16'h04F7;    16'd55249: out <= 16'h059B;    16'd55250: out <= 16'h0244;    16'd55251: out <= 16'hFC33;
    16'd55252: out <= 16'hFE37;    16'd55253: out <= 16'h01FF;    16'd55254: out <= 16'hF416;    16'd55255: out <= 16'h01CD;
    16'd55256: out <= 16'hFE3D;    16'd55257: out <= 16'h0323;    16'd55258: out <= 16'hFFC2;    16'd55259: out <= 16'hFE5D;
    16'd55260: out <= 16'hF9DC;    16'd55261: out <= 16'h085B;    16'd55262: out <= 16'h0580;    16'd55263: out <= 16'hF7FD;
    16'd55264: out <= 16'hFFDE;    16'd55265: out <= 16'h0177;    16'd55266: out <= 16'h03B9;    16'd55267: out <= 16'h038E;
    16'd55268: out <= 16'hFDAF;    16'd55269: out <= 16'h016C;    16'd55270: out <= 16'hFBCC;    16'd55271: out <= 16'h03E8;
    16'd55272: out <= 16'hFD8F;    16'd55273: out <= 16'hF864;    16'd55274: out <= 16'h01D8;    16'd55275: out <= 16'hFFA2;
    16'd55276: out <= 16'h00EC;    16'd55277: out <= 16'hFE1E;    16'd55278: out <= 16'h01DD;    16'd55279: out <= 16'hFE4A;
    16'd55280: out <= 16'hFE27;    16'd55281: out <= 16'hFE56;    16'd55282: out <= 16'h0635;    16'd55283: out <= 16'h063D;
    16'd55284: out <= 16'hFFFB;    16'd55285: out <= 16'hFA24;    16'd55286: out <= 16'hFEFB;    16'd55287: out <= 16'h0286;
    16'd55288: out <= 16'hFCAD;    16'd55289: out <= 16'h0288;    16'd55290: out <= 16'h001F;    16'd55291: out <= 16'h00C3;
    16'd55292: out <= 16'hF95E;    16'd55293: out <= 16'hFBBB;    16'd55294: out <= 16'h0248;    16'd55295: out <= 16'hFA5D;
    16'd55296: out <= 16'hF990;    16'd55297: out <= 16'h01D7;    16'd55298: out <= 16'h02ED;    16'd55299: out <= 16'h04CF;
    16'd55300: out <= 16'hF906;    16'd55301: out <= 16'hFC2D;    16'd55302: out <= 16'h0223;    16'd55303: out <= 16'h03C2;
    16'd55304: out <= 16'hFA19;    16'd55305: out <= 16'hF632;    16'd55306: out <= 16'h0002;    16'd55307: out <= 16'h0159;
    16'd55308: out <= 16'h02C1;    16'd55309: out <= 16'h0078;    16'd55310: out <= 16'hFB23;    16'd55311: out <= 16'h0042;
    16'd55312: out <= 16'h0333;    16'd55313: out <= 16'h0291;    16'd55314: out <= 16'hFF0A;    16'd55315: out <= 16'h0262;
    16'd55316: out <= 16'h0086;    16'd55317: out <= 16'hFC4A;    16'd55318: out <= 16'h03D7;    16'd55319: out <= 16'hFF22;
    16'd55320: out <= 16'h0422;    16'd55321: out <= 16'hFCDE;    16'd55322: out <= 16'hF7DB;    16'd55323: out <= 16'h073C;
    16'd55324: out <= 16'hFE1D;    16'd55325: out <= 16'h006A;    16'd55326: out <= 16'h0551;    16'd55327: out <= 16'hFD70;
    16'd55328: out <= 16'h0098;    16'd55329: out <= 16'h0A6A;    16'd55330: out <= 16'h0087;    16'd55331: out <= 16'h037C;
    16'd55332: out <= 16'h00C9;    16'd55333: out <= 16'hFDF1;    16'd55334: out <= 16'hFDC0;    16'd55335: out <= 16'h0488;
    16'd55336: out <= 16'hFC66;    16'd55337: out <= 16'hFB59;    16'd55338: out <= 16'hFEA3;    16'd55339: out <= 16'hFBAD;
    16'd55340: out <= 16'hFF98;    16'd55341: out <= 16'h07A4;    16'd55342: out <= 16'h034D;    16'd55343: out <= 16'h0023;
    16'd55344: out <= 16'h02A3;    16'd55345: out <= 16'hFF71;    16'd55346: out <= 16'h0332;    16'd55347: out <= 16'h0B0B;
    16'd55348: out <= 16'h05B1;    16'd55349: out <= 16'h00BE;    16'd55350: out <= 16'h032D;    16'd55351: out <= 16'h038D;
    16'd55352: out <= 16'hFA8B;    16'd55353: out <= 16'h01AC;    16'd55354: out <= 16'h0719;    16'd55355: out <= 16'h07A5;
    16'd55356: out <= 16'hFDA3;    16'd55357: out <= 16'h00F2;    16'd55358: out <= 16'h0258;    16'd55359: out <= 16'h065D;
    16'd55360: out <= 16'h02C8;    16'd55361: out <= 16'h062A;    16'd55362: out <= 16'h070C;    16'd55363: out <= 16'h06D1;
    16'd55364: out <= 16'h021C;    16'd55365: out <= 16'h0384;    16'd55366: out <= 16'h0390;    16'd55367: out <= 16'h03F9;
    16'd55368: out <= 16'h07D4;    16'd55369: out <= 16'h08C4;    16'd55370: out <= 16'hFDC0;    16'd55371: out <= 16'h0316;
    16'd55372: out <= 16'h0431;    16'd55373: out <= 16'h016E;    16'd55374: out <= 16'h0430;    16'd55375: out <= 16'h03BD;
    16'd55376: out <= 16'h0442;    16'd55377: out <= 16'h0BD0;    16'd55378: out <= 16'h0854;    16'd55379: out <= 16'h0529;
    16'd55380: out <= 16'h0646;    16'd55381: out <= 16'h0AA9;    16'd55382: out <= 16'hFFFE;    16'd55383: out <= 16'h029B;
    16'd55384: out <= 16'h0A1C;    16'd55385: out <= 16'h01E3;    16'd55386: out <= 16'h058D;    16'd55387: out <= 16'hFE65;
    16'd55388: out <= 16'h06A1;    16'd55389: out <= 16'h01D1;    16'd55390: out <= 16'h0B78;    16'd55391: out <= 16'h0123;
    16'd55392: out <= 16'hFFE6;    16'd55393: out <= 16'hFCC2;    16'd55394: out <= 16'h00ED;    16'd55395: out <= 16'h023A;
    16'd55396: out <= 16'h07F8;    16'd55397: out <= 16'hFF4F;    16'd55398: out <= 16'h0737;    16'd55399: out <= 16'h099D;
    16'd55400: out <= 16'h0681;    16'd55401: out <= 16'h0008;    16'd55402: out <= 16'h0161;    16'd55403: out <= 16'h0719;
    16'd55404: out <= 16'h0152;    16'd55405: out <= 16'h0686;    16'd55406: out <= 16'h0510;    16'd55407: out <= 16'h0464;
    16'd55408: out <= 16'hFFE1;    16'd55409: out <= 16'hFF8D;    16'd55410: out <= 16'h015E;    16'd55411: out <= 16'h0A0B;
    16'd55412: out <= 16'h020C;    16'd55413: out <= 16'h093B;    16'd55414: out <= 16'h0628;    16'd55415: out <= 16'h0A5D;
    16'd55416: out <= 16'h0603;    16'd55417: out <= 16'h044B;    16'd55418: out <= 16'h01FB;    16'd55419: out <= 16'h034B;
    16'd55420: out <= 16'hFFA2;    16'd55421: out <= 16'h0084;    16'd55422: out <= 16'h03FB;    16'd55423: out <= 16'h02E7;
    16'd55424: out <= 16'h002D;    16'd55425: out <= 16'h00E0;    16'd55426: out <= 16'h0438;    16'd55427: out <= 16'h00E1;
    16'd55428: out <= 16'h02DC;    16'd55429: out <= 16'h0049;    16'd55430: out <= 16'h07AA;    16'd55431: out <= 16'hFE25;
    16'd55432: out <= 16'hFEFF;    16'd55433: out <= 16'h0285;    16'd55434: out <= 16'h081B;    16'd55435: out <= 16'hFE36;
    16'd55436: out <= 16'h0249;    16'd55437: out <= 16'h071D;    16'd55438: out <= 16'h032F;    16'd55439: out <= 16'h080A;
    16'd55440: out <= 16'h0876;    16'd55441: out <= 16'h031B;    16'd55442: out <= 16'h03DF;    16'd55443: out <= 16'h01E0;
    16'd55444: out <= 16'h08B0;    16'd55445: out <= 16'h03D4;    16'd55446: out <= 16'h06BB;    16'd55447: out <= 16'h0582;
    16'd55448: out <= 16'h021F;    16'd55449: out <= 16'h02B3;    16'd55450: out <= 16'h03D6;    16'd55451: out <= 16'h005D;
    16'd55452: out <= 16'h09B3;    16'd55453: out <= 16'h0A3C;    16'd55454: out <= 16'h0639;    16'd55455: out <= 16'h00F5;
    16'd55456: out <= 16'h0658;    16'd55457: out <= 16'h0921;    16'd55458: out <= 16'h06D6;    16'd55459: out <= 16'h059C;
    16'd55460: out <= 16'h04F0;    16'd55461: out <= 16'h05FE;    16'd55462: out <= 16'h045F;    16'd55463: out <= 16'hFC67;
    16'd55464: out <= 16'h08F8;    16'd55465: out <= 16'h0707;    16'd55466: out <= 16'h071A;    16'd55467: out <= 16'h02A7;
    16'd55468: out <= 16'h02D7;    16'd55469: out <= 16'hFCBD;    16'd55470: out <= 16'hFD88;    16'd55471: out <= 16'h08FD;
    16'd55472: out <= 16'h0391;    16'd55473: out <= 16'h02AE;    16'd55474: out <= 16'h0537;    16'd55475: out <= 16'h004A;
    16'd55476: out <= 16'h04C9;    16'd55477: out <= 16'h0243;    16'd55478: out <= 16'h08AE;    16'd55479: out <= 16'h04F7;
    16'd55480: out <= 16'h0105;    16'd55481: out <= 16'h03F9;    16'd55482: out <= 16'h05D9;    16'd55483: out <= 16'h065B;
    16'd55484: out <= 16'h05A2;    16'd55485: out <= 16'h03B1;    16'd55486: out <= 16'h05D0;    16'd55487: out <= 16'h03D2;
    16'd55488: out <= 16'h0601;    16'd55489: out <= 16'h06EC;    16'd55490: out <= 16'h0687;    16'd55491: out <= 16'hFDF9;
    16'd55492: out <= 16'hF784;    16'd55493: out <= 16'h02A6;    16'd55494: out <= 16'hFA7E;    16'd55495: out <= 16'h02DA;
    16'd55496: out <= 16'h014C;    16'd55497: out <= 16'hFCB0;    16'd55498: out <= 16'h033F;    16'd55499: out <= 16'h0680;
    16'd55500: out <= 16'hFF29;    16'd55501: out <= 16'hF783;    16'd55502: out <= 16'h0371;    16'd55503: out <= 16'hFA99;
    16'd55504: out <= 16'hFFE8;    16'd55505: out <= 16'hFC76;    16'd55506: out <= 16'h00E1;    16'd55507: out <= 16'hFD4D;
    16'd55508: out <= 16'h0161;    16'd55509: out <= 16'hFEA0;    16'd55510: out <= 16'hFE3B;    16'd55511: out <= 16'h0009;
    16'd55512: out <= 16'hF82B;    16'd55513: out <= 16'h0508;    16'd55514: out <= 16'hFF00;    16'd55515: out <= 16'hFE2F;
    16'd55516: out <= 16'h0065;    16'd55517: out <= 16'h04DF;    16'd55518: out <= 16'hFED4;    16'd55519: out <= 16'hFB82;
    16'd55520: out <= 16'h000C;    16'd55521: out <= 16'hF763;    16'd55522: out <= 16'h0586;    16'd55523: out <= 16'hFEEB;
    16'd55524: out <= 16'h003B;    16'd55525: out <= 16'hFF2D;    16'd55526: out <= 16'hF8F4;    16'd55527: out <= 16'hFFB7;
    16'd55528: out <= 16'hFCC1;    16'd55529: out <= 16'hFFA7;    16'd55530: out <= 16'hFA7C;    16'd55531: out <= 16'hFC05;
    16'd55532: out <= 16'h05E7;    16'd55533: out <= 16'h019F;    16'd55534: out <= 16'hF6DB;    16'd55535: out <= 16'hFD32;
    16'd55536: out <= 16'h034A;    16'd55537: out <= 16'hFC23;    16'd55538: out <= 16'hFDC4;    16'd55539: out <= 16'hF958;
    16'd55540: out <= 16'hFFBB;    16'd55541: out <= 16'h0655;    16'd55542: out <= 16'h070C;    16'd55543: out <= 16'h05D1;
    16'd55544: out <= 16'hFD81;    16'd55545: out <= 16'h027F;    16'd55546: out <= 16'h03F0;    16'd55547: out <= 16'hFCFC;
    16'd55548: out <= 16'hFE8A;    16'd55549: out <= 16'hFC88;    16'd55550: out <= 16'h0106;    16'd55551: out <= 16'hF989;
    16'd55552: out <= 16'h02D9;    16'd55553: out <= 16'h035F;    16'd55554: out <= 16'hFF6E;    16'd55555: out <= 16'hFD7C;
    16'd55556: out <= 16'h0342;    16'd55557: out <= 16'h0562;    16'd55558: out <= 16'hFAB7;    16'd55559: out <= 16'hFD9B;
    16'd55560: out <= 16'h0113;    16'd55561: out <= 16'h0280;    16'd55562: out <= 16'h00CD;    16'd55563: out <= 16'hFE6D;
    16'd55564: out <= 16'hFA20;    16'd55565: out <= 16'h0327;    16'd55566: out <= 16'hFF5A;    16'd55567: out <= 16'h0047;
    16'd55568: out <= 16'h03B8;    16'd55569: out <= 16'hFBFF;    16'd55570: out <= 16'hFDDB;    16'd55571: out <= 16'hFBCD;
    16'd55572: out <= 16'hFE4C;    16'd55573: out <= 16'h050D;    16'd55574: out <= 16'hFEDA;    16'd55575: out <= 16'hFADF;
    16'd55576: out <= 16'hFE39;    16'd55577: out <= 16'hFC93;    16'd55578: out <= 16'h002D;    16'd55579: out <= 16'h007C;
    16'd55580: out <= 16'hFF81;    16'd55581: out <= 16'hFBFF;    16'd55582: out <= 16'hFDDD;    16'd55583: out <= 16'hFE93;
    16'd55584: out <= 16'h00A5;    16'd55585: out <= 16'hFD7A;    16'd55586: out <= 16'hF948;    16'd55587: out <= 16'h01D9;
    16'd55588: out <= 16'h04A0;    16'd55589: out <= 16'h0268;    16'd55590: out <= 16'hFB3F;    16'd55591: out <= 16'hFD23;
    16'd55592: out <= 16'hFC6E;    16'd55593: out <= 16'hFBD8;    16'd55594: out <= 16'h0184;    16'd55595: out <= 16'hFBF5;
    16'd55596: out <= 16'h0374;    16'd55597: out <= 16'h0323;    16'd55598: out <= 16'h026E;    16'd55599: out <= 16'hFF39;
    16'd55600: out <= 16'h0147;    16'd55601: out <= 16'h0414;    16'd55602: out <= 16'h0576;    16'd55603: out <= 16'hFC3C;
    16'd55604: out <= 16'h03F2;    16'd55605: out <= 16'h0736;    16'd55606: out <= 16'h036F;    16'd55607: out <= 16'h081B;
    16'd55608: out <= 16'h06A7;    16'd55609: out <= 16'h02DC;    16'd55610: out <= 16'h0AAF;    16'd55611: out <= 16'h0696;
    16'd55612: out <= 16'h08E9;    16'd55613: out <= 16'h0284;    16'd55614: out <= 16'h07B4;    16'd55615: out <= 16'h061A;
    16'd55616: out <= 16'h0226;    16'd55617: out <= 16'h0F9C;    16'd55618: out <= 16'h0165;    16'd55619: out <= 16'h0732;
    16'd55620: out <= 16'h097A;    16'd55621: out <= 16'h0737;    16'd55622: out <= 16'hFC36;    16'd55623: out <= 16'h0899;
    16'd55624: out <= 16'hFFA5;    16'd55625: out <= 16'h054F;    16'd55626: out <= 16'h0A1F;    16'd55627: out <= 16'h08AD;
    16'd55628: out <= 16'h05B0;    16'd55629: out <= 16'h0152;    16'd55630: out <= 16'hFD2F;    16'd55631: out <= 16'h0459;
    16'd55632: out <= 16'h0415;    16'd55633: out <= 16'h0546;    16'd55634: out <= 16'h09AB;    16'd55635: out <= 16'h03E5;
    16'd55636: out <= 16'h01C7;    16'd55637: out <= 16'hFEF8;    16'd55638: out <= 16'h01FE;    16'd55639: out <= 16'hFCDD;
    16'd55640: out <= 16'h0256;    16'd55641: out <= 16'h06D0;    16'd55642: out <= 16'h04FC;    16'd55643: out <= 16'h0344;
    16'd55644: out <= 16'h0327;    16'd55645: out <= 16'h038D;    16'd55646: out <= 16'h07B9;    16'd55647: out <= 16'h0641;
    16'd55648: out <= 16'hFFCD;    16'd55649: out <= 16'h038E;    16'd55650: out <= 16'h0508;    16'd55651: out <= 16'h058E;
    16'd55652: out <= 16'hFE68;    16'd55653: out <= 16'h01D1;    16'd55654: out <= 16'h089A;    16'd55655: out <= 16'h05EF;
    16'd55656: out <= 16'h05BD;    16'd55657: out <= 16'h03CB;    16'd55658: out <= 16'h007D;    16'd55659: out <= 16'h0102;
    16'd55660: out <= 16'h089B;    16'd55661: out <= 16'h07FB;    16'd55662: out <= 16'hFCE0;    16'd55663: out <= 16'h06A0;
    16'd55664: out <= 16'h09BD;    16'd55665: out <= 16'h0894;    16'd55666: out <= 16'h03C8;    16'd55667: out <= 16'h0495;
    16'd55668: out <= 16'h05A4;    16'd55669: out <= 16'h078C;    16'd55670: out <= 16'h03DF;    16'd55671: out <= 16'hFF8A;
    16'd55672: out <= 16'h0138;    16'd55673: out <= 16'h0640;    16'd55674: out <= 16'h07BF;    16'd55675: out <= 16'h03B8;
    16'd55676: out <= 16'h0AED;    16'd55677: out <= 16'h005B;    16'd55678: out <= 16'h0748;    16'd55679: out <= 16'h0566;
    16'd55680: out <= 16'h0304;    16'd55681: out <= 16'hFF4E;    16'd55682: out <= 16'h04ED;    16'd55683: out <= 16'h084E;
    16'd55684: out <= 16'h0BA4;    16'd55685: out <= 16'h0217;    16'd55686: out <= 16'h043A;    16'd55687: out <= 16'h05D7;
    16'd55688: out <= 16'h069E;    16'd55689: out <= 16'h0273;    16'd55690: out <= 16'hFE87;    16'd55691: out <= 16'h016A;
    16'd55692: out <= 16'hFCDF;    16'd55693: out <= 16'h015F;    16'd55694: out <= 16'h02CB;    16'd55695: out <= 16'h02CB;
    16'd55696: out <= 16'hFE36;    16'd55697: out <= 16'h0067;    16'd55698: out <= 16'h0467;    16'd55699: out <= 16'hFF43;
    16'd55700: out <= 16'h0200;    16'd55701: out <= 16'h039B;    16'd55702: out <= 16'hFBEC;    16'd55703: out <= 16'h0397;
    16'd55704: out <= 16'h04EC;    16'd55705: out <= 16'h055D;    16'd55706: out <= 16'h0B7D;    16'd55707: out <= 16'h0231;
    16'd55708: out <= 16'h0124;    16'd55709: out <= 16'h015C;    16'd55710: out <= 16'h085E;    16'd55711: out <= 16'h0538;
    16'd55712: out <= 16'h06FA;    16'd55713: out <= 16'h019C;    16'd55714: out <= 16'h0333;    16'd55715: out <= 16'h0242;
    16'd55716: out <= 16'h055B;    16'd55717: out <= 16'h022C;    16'd55718: out <= 16'h06FE;    16'd55719: out <= 16'h05A9;
    16'd55720: out <= 16'h0999;    16'd55721: out <= 16'h08E5;    16'd55722: out <= 16'h0E1E;    16'd55723: out <= 16'h0B0D;
    16'd55724: out <= 16'h0150;    16'd55725: out <= 16'hFE1B;    16'd55726: out <= 16'h074B;    16'd55727: out <= 16'h039A;
    16'd55728: out <= 16'h08A1;    16'd55729: out <= 16'h011F;    16'd55730: out <= 16'hFD73;    16'd55731: out <= 16'hFF7F;
    16'd55732: out <= 16'h047A;    16'd55733: out <= 16'h0896;    16'd55734: out <= 16'h0299;    16'd55735: out <= 16'h07B7;
    16'd55736: out <= 16'h00B6;    16'd55737: out <= 16'h01F6;    16'd55738: out <= 16'h039D;    16'd55739: out <= 16'h0663;
    16'd55740: out <= 16'h0C01;    16'd55741: out <= 16'h08F8;    16'd55742: out <= 16'h034C;    16'd55743: out <= 16'h0577;
    16'd55744: out <= 16'h0514;    16'd55745: out <= 16'h0859;    16'd55746: out <= 16'h0989;    16'd55747: out <= 16'hFB9C;
    16'd55748: out <= 16'hFF03;    16'd55749: out <= 16'h0361;    16'd55750: out <= 16'hFE87;    16'd55751: out <= 16'hFE1E;
    16'd55752: out <= 16'hFA25;    16'd55753: out <= 16'h030E;    16'd55754: out <= 16'h02C8;    16'd55755: out <= 16'h0687;
    16'd55756: out <= 16'h00E3;    16'd55757: out <= 16'hFF2F;    16'd55758: out <= 16'h0313;    16'd55759: out <= 16'h0053;
    16'd55760: out <= 16'h0514;    16'd55761: out <= 16'hFD9F;    16'd55762: out <= 16'h05AE;    16'd55763: out <= 16'hFA55;
    16'd55764: out <= 16'hFAB4;    16'd55765: out <= 16'hFE05;    16'd55766: out <= 16'h039E;    16'd55767: out <= 16'h0710;
    16'd55768: out <= 16'hFDF0;    16'd55769: out <= 16'h00FF;    16'd55770: out <= 16'h0182;    16'd55771: out <= 16'hFD4B;
    16'd55772: out <= 16'h0117;    16'd55773: out <= 16'hFE42;    16'd55774: out <= 16'hFCAF;    16'd55775: out <= 16'hFBD8;
    16'd55776: out <= 16'hFE78;    16'd55777: out <= 16'hFC95;    16'd55778: out <= 16'hFA87;    16'd55779: out <= 16'hFEEF;
    16'd55780: out <= 16'hF97B;    16'd55781: out <= 16'h06BB;    16'd55782: out <= 16'h02C8;    16'd55783: out <= 16'h013E;
    16'd55784: out <= 16'h0A9A;    16'd55785: out <= 16'h06DC;    16'd55786: out <= 16'h0088;    16'd55787: out <= 16'h0462;
    16'd55788: out <= 16'h03AE;    16'd55789: out <= 16'h0339;    16'd55790: out <= 16'hFD1F;    16'd55791: out <= 16'hFFAD;
    16'd55792: out <= 16'hF9B7;    16'd55793: out <= 16'h02CC;    16'd55794: out <= 16'h04C2;    16'd55795: out <= 16'hFE9F;
    16'd55796: out <= 16'h0183;    16'd55797: out <= 16'hFFA8;    16'd55798: out <= 16'hFE70;    16'd55799: out <= 16'hFD83;
    16'd55800: out <= 16'h031D;    16'd55801: out <= 16'hFC40;    16'd55802: out <= 16'hFC74;    16'd55803: out <= 16'hFFC3;
    16'd55804: out <= 16'h050B;    16'd55805: out <= 16'h00D9;    16'd55806: out <= 16'hF918;    16'd55807: out <= 16'h0144;
    16'd55808: out <= 16'hFFA3;    16'd55809: out <= 16'h01DE;    16'd55810: out <= 16'h03DB;    16'd55811: out <= 16'hFEDE;
    16'd55812: out <= 16'hFFBD;    16'd55813: out <= 16'hF5CF;    16'd55814: out <= 16'h032B;    16'd55815: out <= 16'h030B;
    16'd55816: out <= 16'hFFF8;    16'd55817: out <= 16'hFBE4;    16'd55818: out <= 16'hFD67;    16'd55819: out <= 16'h011F;
    16'd55820: out <= 16'hFF75;    16'd55821: out <= 16'hFD23;    16'd55822: out <= 16'h05E5;    16'd55823: out <= 16'h0436;
    16'd55824: out <= 16'hFC57;    16'd55825: out <= 16'h031D;    16'd55826: out <= 16'hFDF1;    16'd55827: out <= 16'hFF15;
    16'd55828: out <= 16'hFDF7;    16'd55829: out <= 16'h05E1;    16'd55830: out <= 16'h002F;    16'd55831: out <= 16'hFF17;
    16'd55832: out <= 16'h0570;    16'd55833: out <= 16'h0130;    16'd55834: out <= 16'h029B;    16'd55835: out <= 16'hFF0D;
    16'd55836: out <= 16'h00F8;    16'd55837: out <= 16'h006D;    16'd55838: out <= 16'hFCDC;    16'd55839: out <= 16'hFF0C;
    16'd55840: out <= 16'h00F8;    16'd55841: out <= 16'h0047;    16'd55842: out <= 16'h0157;    16'd55843: out <= 16'hF7D9;
    16'd55844: out <= 16'hFE2E;    16'd55845: out <= 16'h04AE;    16'd55846: out <= 16'h01ED;    16'd55847: out <= 16'h01F5;
    16'd55848: out <= 16'h01B9;    16'd55849: out <= 16'h003E;    16'd55850: out <= 16'h03A6;    16'd55851: out <= 16'h029A;
    16'd55852: out <= 16'h0090;    16'd55853: out <= 16'h0165;    16'd55854: out <= 16'h06B4;    16'd55855: out <= 16'hFDB5;
    16'd55856: out <= 16'h015D;    16'd55857: out <= 16'hFF04;    16'd55858: out <= 16'h03D9;    16'd55859: out <= 16'h0B27;
    16'd55860: out <= 16'hFFA9;    16'd55861: out <= 16'h0859;    16'd55862: out <= 16'h0231;    16'd55863: out <= 16'hFEFF;
    16'd55864: out <= 16'h08E8;    16'd55865: out <= 16'h0600;    16'd55866: out <= 16'h0342;    16'd55867: out <= 16'h00AB;
    16'd55868: out <= 16'h02A7;    16'd55869: out <= 16'h0097;    16'd55870: out <= 16'h04CA;    16'd55871: out <= 16'h059C;
    16'd55872: out <= 16'hFD60;    16'd55873: out <= 16'h0021;    16'd55874: out <= 16'hFE47;    16'd55875: out <= 16'h0184;
    16'd55876: out <= 16'h086C;    16'd55877: out <= 16'h0E55;    16'd55878: out <= 16'h046C;    16'd55879: out <= 16'h00A3;
    16'd55880: out <= 16'h02C7;    16'd55881: out <= 16'h06D6;    16'd55882: out <= 16'h03D6;    16'd55883: out <= 16'h05B8;
    16'd55884: out <= 16'h0C8C;    16'd55885: out <= 16'h03C0;    16'd55886: out <= 16'h051B;    16'd55887: out <= 16'hFECF;
    16'd55888: out <= 16'h006C;    16'd55889: out <= 16'h0A1A;    16'd55890: out <= 16'h0295;    16'd55891: out <= 16'hFFE5;
    16'd55892: out <= 16'h0253;    16'd55893: out <= 16'h03BD;    16'd55894: out <= 16'h0604;    16'd55895: out <= 16'h02BD;
    16'd55896: out <= 16'h02F7;    16'd55897: out <= 16'hFF2B;    16'd55898: out <= 16'h00A2;    16'd55899: out <= 16'h004C;
    16'd55900: out <= 16'h01CB;    16'd55901: out <= 16'h0455;    16'd55902: out <= 16'h04AE;    16'd55903: out <= 16'h0303;
    16'd55904: out <= 16'h0640;    16'd55905: out <= 16'h0355;    16'd55906: out <= 16'h0835;    16'd55907: out <= 16'h012B;
    16'd55908: out <= 16'h0039;    16'd55909: out <= 16'h04A5;    16'd55910: out <= 16'h02E3;    16'd55911: out <= 16'h0303;
    16'd55912: out <= 16'h041C;    16'd55913: out <= 16'hFFFB;    16'd55914: out <= 16'h08EC;    16'd55915: out <= 16'h0DD2;
    16'd55916: out <= 16'h01B8;    16'd55917: out <= 16'h0150;    16'd55918: out <= 16'h03AD;    16'd55919: out <= 16'h0798;
    16'd55920: out <= 16'hFD3D;    16'd55921: out <= 16'h031E;    16'd55922: out <= 16'h0902;    16'd55923: out <= 16'h0580;
    16'd55924: out <= 16'h0608;    16'd55925: out <= 16'h084B;    16'd55926: out <= 16'h073B;    16'd55927: out <= 16'h0062;
    16'd55928: out <= 16'h0A39;    16'd55929: out <= 16'hFB9E;    16'd55930: out <= 16'h0088;    16'd55931: out <= 16'h0683;
    16'd55932: out <= 16'h06CD;    16'd55933: out <= 16'hFEFC;    16'd55934: out <= 16'h06AD;    16'd55935: out <= 16'h04C9;
    16'd55936: out <= 16'h0492;    16'd55937: out <= 16'h06ED;    16'd55938: out <= 16'h0088;    16'd55939: out <= 16'h042C;
    16'd55940: out <= 16'h026A;    16'd55941: out <= 16'h03E9;    16'd55942: out <= 16'h0511;    16'd55943: out <= 16'h09A7;
    16'd55944: out <= 16'h07B1;    16'd55945: out <= 16'h005E;    16'd55946: out <= 16'h004A;    16'd55947: out <= 16'h0783;
    16'd55948: out <= 16'h0BE8;    16'd55949: out <= 16'h07B7;    16'd55950: out <= 16'h0615;    16'd55951: out <= 16'hFDC5;
    16'd55952: out <= 16'hFC3C;    16'd55953: out <= 16'h063A;    16'd55954: out <= 16'h0040;    16'd55955: out <= 16'h049F;
    16'd55956: out <= 16'h05C2;    16'd55957: out <= 16'h0314;    16'd55958: out <= 16'h01ED;    16'd55959: out <= 16'hFC50;
    16'd55960: out <= 16'h091F;    16'd55961: out <= 16'h0353;    16'd55962: out <= 16'h0583;    16'd55963: out <= 16'h019F;
    16'd55964: out <= 16'hFF00;    16'd55965: out <= 16'h04EF;    16'd55966: out <= 16'hFF2D;    16'd55967: out <= 16'h05FC;
    16'd55968: out <= 16'hFE45;    16'd55969: out <= 16'h051E;    16'd55970: out <= 16'h0B5E;    16'd55971: out <= 16'h0165;
    16'd55972: out <= 16'h06BD;    16'd55973: out <= 16'h03DF;    16'd55974: out <= 16'h0A2C;    16'd55975: out <= 16'h0016;
    16'd55976: out <= 16'h0095;    16'd55977: out <= 16'h040E;    16'd55978: out <= 16'h06FA;    16'd55979: out <= 16'h0462;
    16'd55980: out <= 16'h005E;    16'd55981: out <= 16'h04A0;    16'd55982: out <= 16'h076A;    16'd55983: out <= 16'h0695;
    16'd55984: out <= 16'h03DC;    16'd55985: out <= 16'h0756;    16'd55986: out <= 16'hF927;    16'd55987: out <= 16'h05A5;
    16'd55988: out <= 16'h044B;    16'd55989: out <= 16'hFE2D;    16'd55990: out <= 16'h05A2;    16'd55991: out <= 16'h0150;
    16'd55992: out <= 16'h044A;    16'd55993: out <= 16'h0891;    16'd55994: out <= 16'hFE4D;    16'd55995: out <= 16'h0231;
    16'd55996: out <= 16'h0557;    16'd55997: out <= 16'h0596;    16'd55998: out <= 16'h0B80;    16'd55999: out <= 16'hFBDD;
    16'd56000: out <= 16'h0457;    16'd56001: out <= 16'h0499;    16'd56002: out <= 16'h08E5;    16'd56003: out <= 16'hF883;
    16'd56004: out <= 16'h0232;    16'd56005: out <= 16'hF74F;    16'd56006: out <= 16'h05AC;    16'd56007: out <= 16'hFE1B;
    16'd56008: out <= 16'h03A6;    16'd56009: out <= 16'hFFFA;    16'd56010: out <= 16'h02A7;    16'd56011: out <= 16'h0174;
    16'd56012: out <= 16'hF9FA;    16'd56013: out <= 16'h091E;    16'd56014: out <= 16'h0356;    16'd56015: out <= 16'h0664;
    16'd56016: out <= 16'h0237;    16'd56017: out <= 16'hFB5B;    16'd56018: out <= 16'h0151;    16'd56019: out <= 16'h018E;
    16'd56020: out <= 16'h033C;    16'd56021: out <= 16'hFDF9;    16'd56022: out <= 16'h0597;    16'd56023: out <= 16'h064A;
    16'd56024: out <= 16'h051D;    16'd56025: out <= 16'hFC67;    16'd56026: out <= 16'h02DE;    16'd56027: out <= 16'hFF5C;
    16'd56028: out <= 16'hFBA2;    16'd56029: out <= 16'h004D;    16'd56030: out <= 16'h010A;    16'd56031: out <= 16'h0670;
    16'd56032: out <= 16'h0668;    16'd56033: out <= 16'h0228;    16'd56034: out <= 16'h078F;    16'd56035: out <= 16'h0432;
    16'd56036: out <= 16'hFD45;    16'd56037: out <= 16'h00DD;    16'd56038: out <= 16'hFE01;    16'd56039: out <= 16'h0145;
    16'd56040: out <= 16'hFADB;    16'd56041: out <= 16'h07B3;    16'd56042: out <= 16'hFF29;    16'd56043: out <= 16'hFDB9;
    16'd56044: out <= 16'hF81B;    16'd56045: out <= 16'hFDA1;    16'd56046: out <= 16'hFF5F;    16'd56047: out <= 16'h0401;
    16'd56048: out <= 16'h040A;    16'd56049: out <= 16'h00CF;    16'd56050: out <= 16'hFECF;    16'd56051: out <= 16'h027D;
    16'd56052: out <= 16'hFABE;    16'd56053: out <= 16'h0723;    16'd56054: out <= 16'hF8F1;    16'd56055: out <= 16'h0209;
    16'd56056: out <= 16'hFCE9;    16'd56057: out <= 16'h0405;    16'd56058: out <= 16'h00F3;    16'd56059: out <= 16'h01B5;
    16'd56060: out <= 16'hFC41;    16'd56061: out <= 16'h07B2;    16'd56062: out <= 16'hFBC0;    16'd56063: out <= 16'h0765;
    16'd56064: out <= 16'hFA1E;    16'd56065: out <= 16'h0003;    16'd56066: out <= 16'h023B;    16'd56067: out <= 16'hFDAD;
    16'd56068: out <= 16'h0105;    16'd56069: out <= 16'h05E5;    16'd56070: out <= 16'h02E1;    16'd56071: out <= 16'h0024;
    16'd56072: out <= 16'h009B;    16'd56073: out <= 16'hFACA;    16'd56074: out <= 16'hFD7C;    16'd56075: out <= 16'h07C1;
    16'd56076: out <= 16'h0217;    16'd56077: out <= 16'hFC39;    16'd56078: out <= 16'hFD16;    16'd56079: out <= 16'hFEB9;
    16'd56080: out <= 16'hFB43;    16'd56081: out <= 16'h04C3;    16'd56082: out <= 16'h0128;    16'd56083: out <= 16'hFF28;
    16'd56084: out <= 16'h02A1;    16'd56085: out <= 16'h01FA;    16'd56086: out <= 16'hFC0D;    16'd56087: out <= 16'h02B6;
    16'd56088: out <= 16'hFE09;    16'd56089: out <= 16'hFCA0;    16'd56090: out <= 16'hFA34;    16'd56091: out <= 16'h0296;
    16'd56092: out <= 16'h0095;    16'd56093: out <= 16'h0122;    16'd56094: out <= 16'h00EA;    16'd56095: out <= 16'h0098;
    16'd56096: out <= 16'hF4B0;    16'd56097: out <= 16'hFF3F;    16'd56098: out <= 16'h06BD;    16'd56099: out <= 16'hFC66;
    16'd56100: out <= 16'hFC68;    16'd56101: out <= 16'hFD5D;    16'd56102: out <= 16'h04DC;    16'd56103: out <= 16'h0089;
    16'd56104: out <= 16'h004A;    16'd56105: out <= 16'hFAD7;    16'd56106: out <= 16'hFBE6;    16'd56107: out <= 16'h024C;
    16'd56108: out <= 16'h01EA;    16'd56109: out <= 16'hFBFA;    16'd56110: out <= 16'h008C;    16'd56111: out <= 16'h03F2;
    16'd56112: out <= 16'h0375;    16'd56113: out <= 16'h05BA;    16'd56114: out <= 16'h0599;    16'd56115: out <= 16'h0005;
    16'd56116: out <= 16'hFF86;    16'd56117: out <= 16'h0412;    16'd56118: out <= 16'h0244;    16'd56119: out <= 16'h05EB;
    16'd56120: out <= 16'h01A8;    16'd56121: out <= 16'h031F;    16'd56122: out <= 16'h02C5;    16'd56123: out <= 16'h022D;
    16'd56124: out <= 16'h0034;    16'd56125: out <= 16'h00CC;    16'd56126: out <= 16'hFCB1;    16'd56127: out <= 16'h067C;
    16'd56128: out <= 16'h0704;    16'd56129: out <= 16'h0226;    16'd56130: out <= 16'h0213;    16'd56131: out <= 16'h0575;
    16'd56132: out <= 16'h0136;    16'd56133: out <= 16'h0626;    16'd56134: out <= 16'hF61D;    16'd56135: out <= 16'h0390;
    16'd56136: out <= 16'hFE1A;    16'd56137: out <= 16'hFAD6;    16'd56138: out <= 16'h058A;    16'd56139: out <= 16'hFF7B;
    16'd56140: out <= 16'hFCA1;    16'd56141: out <= 16'h060A;    16'd56142: out <= 16'h005E;    16'd56143: out <= 16'hFDC7;
    16'd56144: out <= 16'h0462;    16'd56145: out <= 16'h0594;    16'd56146: out <= 16'hFE2E;    16'd56147: out <= 16'h00CD;
    16'd56148: out <= 16'h005B;    16'd56149: out <= 16'h0049;    16'd56150: out <= 16'h021E;    16'd56151: out <= 16'h029E;
    16'd56152: out <= 16'h0436;    16'd56153: out <= 16'h03BB;    16'd56154: out <= 16'h0AA8;    16'd56155: out <= 16'h01C2;
    16'd56156: out <= 16'h09AF;    16'd56157: out <= 16'hFF07;    16'd56158: out <= 16'h0408;    16'd56159: out <= 16'h0017;
    16'd56160: out <= 16'h0217;    16'd56161: out <= 16'h068F;    16'd56162: out <= 16'h032C;    16'd56163: out <= 16'h088A;
    16'd56164: out <= 16'h029F;    16'd56165: out <= 16'h0443;    16'd56166: out <= 16'h0130;    16'd56167: out <= 16'h0589;
    16'd56168: out <= 16'h01FC;    16'd56169: out <= 16'h037C;    16'd56170: out <= 16'h034A;    16'd56171: out <= 16'h0670;
    16'd56172: out <= 16'h0959;    16'd56173: out <= 16'hFF57;    16'd56174: out <= 16'h078B;    16'd56175: out <= 16'h080E;
    16'd56176: out <= 16'h0649;    16'd56177: out <= 16'h038D;    16'd56178: out <= 16'hFE77;    16'd56179: out <= 16'h073D;
    16'd56180: out <= 16'h06E9;    16'd56181: out <= 16'hFD4E;    16'd56182: out <= 16'h041A;    16'd56183: out <= 16'h0E01;
    16'd56184: out <= 16'h0655;    16'd56185: out <= 16'h0D6C;    16'd56186: out <= 16'h0722;    16'd56187: out <= 16'h0643;
    16'd56188: out <= 16'h07FA;    16'd56189: out <= 16'h0129;    16'd56190: out <= 16'h0071;    16'd56191: out <= 16'h080F;
    16'd56192: out <= 16'h0BBA;    16'd56193: out <= 16'h012F;    16'd56194: out <= 16'hFC34;    16'd56195: out <= 16'h0166;
    16'd56196: out <= 16'hFEE7;    16'd56197: out <= 16'h04EA;    16'd56198: out <= 16'h01A4;    16'd56199: out <= 16'h0371;
    16'd56200: out <= 16'hFE3E;    16'd56201: out <= 16'h05B8;    16'd56202: out <= 16'h0475;    16'd56203: out <= 16'h08BB;
    16'd56204: out <= 16'h027A;    16'd56205: out <= 16'hFDBD;    16'd56206: out <= 16'h04CB;    16'd56207: out <= 16'h0803;
    16'd56208: out <= 16'h0C52;    16'd56209: out <= 16'h059C;    16'd56210: out <= 16'h0408;    16'd56211: out <= 16'h068E;
    16'd56212: out <= 16'hFC93;    16'd56213: out <= 16'h01F4;    16'd56214: out <= 16'h07FB;    16'd56215: out <= 16'h0219;
    16'd56216: out <= 16'h0445;    16'd56217: out <= 16'h076A;    16'd56218: out <= 16'h0367;    16'd56219: out <= 16'h0B67;
    16'd56220: out <= 16'hFF88;    16'd56221: out <= 16'hFFDB;    16'd56222: out <= 16'h00F4;    16'd56223: out <= 16'h06D0;
    16'd56224: out <= 16'h0226;    16'd56225: out <= 16'h01BB;    16'd56226: out <= 16'h03F7;    16'd56227: out <= 16'hFC79;
    16'd56228: out <= 16'h0787;    16'd56229: out <= 16'h0003;    16'd56230: out <= 16'hFF18;    16'd56231: out <= 16'h0707;
    16'd56232: out <= 16'h06DF;    16'd56233: out <= 16'hFE68;    16'd56234: out <= 16'h03B3;    16'd56235: out <= 16'h0690;
    16'd56236: out <= 16'h09B9;    16'd56237: out <= 16'h05D9;    16'd56238: out <= 16'h03C9;    16'd56239: out <= 16'h050C;
    16'd56240: out <= 16'h03EA;    16'd56241: out <= 16'h02DB;    16'd56242: out <= 16'h0765;    16'd56243: out <= 16'hFF47;
    16'd56244: out <= 16'h0478;    16'd56245: out <= 16'hFE98;    16'd56246: out <= 16'h065F;    16'd56247: out <= 16'h08C2;
    16'd56248: out <= 16'hFED0;    16'd56249: out <= 16'h0B9C;    16'd56250: out <= 16'h0329;    16'd56251: out <= 16'h010F;
    16'd56252: out <= 16'h0273;    16'd56253: out <= 16'h0888;    16'd56254: out <= 16'h0385;    16'd56255: out <= 16'h09A0;
    16'd56256: out <= 16'hFFDB;    16'd56257: out <= 16'h08D3;    16'd56258: out <= 16'h063A;    16'd56259: out <= 16'h0566;
    16'd56260: out <= 16'hFD13;    16'd56261: out <= 16'h01CC;    16'd56262: out <= 16'h00BD;    16'd56263: out <= 16'hFDCF;
    16'd56264: out <= 16'h0546;    16'd56265: out <= 16'hFD9F;    16'd56266: out <= 16'h0301;    16'd56267: out <= 16'h0263;
    16'd56268: out <= 16'h0101;    16'd56269: out <= 16'hFC34;    16'd56270: out <= 16'h001F;    16'd56271: out <= 16'hFDAE;
    16'd56272: out <= 16'h025F;    16'd56273: out <= 16'h05A8;    16'd56274: out <= 16'h00DF;    16'd56275: out <= 16'h0285;
    16'd56276: out <= 16'h00B7;    16'd56277: out <= 16'h0175;    16'd56278: out <= 16'h0183;    16'd56279: out <= 16'hFDD8;
    16'd56280: out <= 16'h071D;    16'd56281: out <= 16'hFE34;    16'd56282: out <= 16'h0123;    16'd56283: out <= 16'hFF4C;
    16'd56284: out <= 16'hF87D;    16'd56285: out <= 16'hFD60;    16'd56286: out <= 16'hFF03;    16'd56287: out <= 16'hFBC7;
    16'd56288: out <= 16'hFA21;    16'd56289: out <= 16'hFFEC;    16'd56290: out <= 16'h01FC;    16'd56291: out <= 16'h01D2;
    16'd56292: out <= 16'h015B;    16'd56293: out <= 16'hFD15;    16'd56294: out <= 16'hFEDC;    16'd56295: out <= 16'h08FF;
    16'd56296: out <= 16'h021C;    16'd56297: out <= 16'hFE36;    16'd56298: out <= 16'hFC13;    16'd56299: out <= 16'h0520;
    16'd56300: out <= 16'hFEFE;    16'd56301: out <= 16'h0395;    16'd56302: out <= 16'hFCEC;    16'd56303: out <= 16'h00EF;
    16'd56304: out <= 16'hFBE7;    16'd56305: out <= 16'h035A;    16'd56306: out <= 16'h02CD;    16'd56307: out <= 16'hFC1F;
    16'd56308: out <= 16'h05B3;    16'd56309: out <= 16'h01C2;    16'd56310: out <= 16'hFA9E;    16'd56311: out <= 16'h0369;
    16'd56312: out <= 16'hFBA2;    16'd56313: out <= 16'hFE11;    16'd56314: out <= 16'hFF85;    16'd56315: out <= 16'hFACE;
    16'd56316: out <= 16'h0355;    16'd56317: out <= 16'h020D;    16'd56318: out <= 16'h0880;    16'd56319: out <= 16'h00B8;
    16'd56320: out <= 16'hFFB5;    16'd56321: out <= 16'h00E3;    16'd56322: out <= 16'hFB79;    16'd56323: out <= 16'h007D;
    16'd56324: out <= 16'hFD33;    16'd56325: out <= 16'h0090;    16'd56326: out <= 16'hFE6E;    16'd56327: out <= 16'hFD99;
    16'd56328: out <= 16'hFE7E;    16'd56329: out <= 16'hFD86;    16'd56330: out <= 16'hFB92;    16'd56331: out <= 16'h0605;
    16'd56332: out <= 16'hFF9D;    16'd56333: out <= 16'h0458;    16'd56334: out <= 16'hFF4D;    16'd56335: out <= 16'hFBC6;
    16'd56336: out <= 16'h00DC;    16'd56337: out <= 16'h01A4;    16'd56338: out <= 16'hFD06;    16'd56339: out <= 16'h05FC;
    16'd56340: out <= 16'hFF15;    16'd56341: out <= 16'hFA2B;    16'd56342: out <= 16'h0106;    16'd56343: out <= 16'hFA52;
    16'd56344: out <= 16'hFADC;    16'd56345: out <= 16'hFE88;    16'd56346: out <= 16'h00C4;    16'd56347: out <= 16'hFCD7;
    16'd56348: out <= 16'hFD19;    16'd56349: out <= 16'hFCE1;    16'd56350: out <= 16'hFE3A;    16'd56351: out <= 16'hFD05;
    16'd56352: out <= 16'hFC94;    16'd56353: out <= 16'h0303;    16'd56354: out <= 16'h02EF;    16'd56355: out <= 16'hFD17;
    16'd56356: out <= 16'hFEFA;    16'd56357: out <= 16'hF7E6;    16'd56358: out <= 16'h0389;    16'd56359: out <= 16'hFFB4;
    16'd56360: out <= 16'hFCAA;    16'd56361: out <= 16'hFF72;    16'd56362: out <= 16'h020C;    16'd56363: out <= 16'h0028;
    16'd56364: out <= 16'hFE99;    16'd56365: out <= 16'h086C;    16'd56366: out <= 16'h004C;    16'd56367: out <= 16'hFD57;
    16'd56368: out <= 16'h09C0;    16'd56369: out <= 16'h00F2;    16'd56370: out <= 16'h015C;    16'd56371: out <= 16'hFD71;
    16'd56372: out <= 16'hFF02;    16'd56373: out <= 16'hFFA6;    16'd56374: out <= 16'h0443;    16'd56375: out <= 16'h0518;
    16'd56376: out <= 16'h0693;    16'd56377: out <= 16'h0192;    16'd56378: out <= 16'h04EF;    16'd56379: out <= 16'h0B6E;
    16'd56380: out <= 16'h0310;    16'd56381: out <= 16'h079B;    16'd56382: out <= 16'h0324;    16'd56383: out <= 16'h0893;
    16'd56384: out <= 16'h084C;    16'd56385: out <= 16'h0B16;    16'd56386: out <= 16'h0302;    16'd56387: out <= 16'h0762;
    16'd56388: out <= 16'h0855;    16'd56389: out <= 16'h07FE;    16'd56390: out <= 16'h02F0;    16'd56391: out <= 16'h029C;
    16'd56392: out <= 16'hFECF;    16'd56393: out <= 16'h089A;    16'd56394: out <= 16'h003D;    16'd56395: out <= 16'h0CEB;
    16'd56396: out <= 16'h02B3;    16'd56397: out <= 16'h0104;    16'd56398: out <= 16'h03EA;    16'd56399: out <= 16'h039A;
    16'd56400: out <= 16'h0343;    16'd56401: out <= 16'h05BB;    16'd56402: out <= 16'h017A;    16'd56403: out <= 16'h01B5;
    16'd56404: out <= 16'h044D;    16'd56405: out <= 16'h0402;    16'd56406: out <= 16'h06E5;    16'd56407: out <= 16'h05BA;
    16'd56408: out <= 16'h019D;    16'd56409: out <= 16'hFE43;    16'd56410: out <= 16'h0048;    16'd56411: out <= 16'hFEF3;
    16'd56412: out <= 16'h066C;    16'd56413: out <= 16'h00A7;    16'd56414: out <= 16'h0ABD;    16'd56415: out <= 16'h0993;
    16'd56416: out <= 16'hFCF8;    16'd56417: out <= 16'h00E9;    16'd56418: out <= 16'h0181;    16'd56419: out <= 16'hFE9A;
    16'd56420: out <= 16'h05A1;    16'd56421: out <= 16'h07A4;    16'd56422: out <= 16'hFB28;    16'd56423: out <= 16'h0062;
    16'd56424: out <= 16'h05A1;    16'd56425: out <= 16'h0747;    16'd56426: out <= 16'h03D0;    16'd56427: out <= 16'h05F3;
    16'd56428: out <= 16'hFDAC;    16'd56429: out <= 16'hFF8D;    16'd56430: out <= 16'hFBC2;    16'd56431: out <= 16'h0440;
    16'd56432: out <= 16'h03D9;    16'd56433: out <= 16'h00D1;    16'd56434: out <= 16'h0402;    16'd56435: out <= 16'h0794;
    16'd56436: out <= 16'h07EE;    16'd56437: out <= 16'hFEC8;    16'd56438: out <= 16'h027A;    16'd56439: out <= 16'h046A;
    16'd56440: out <= 16'h01AD;    16'd56441: out <= 16'h03CA;    16'd56442: out <= 16'h0626;    16'd56443: out <= 16'h040D;
    16'd56444: out <= 16'h0437;    16'd56445: out <= 16'hFBB7;    16'd56446: out <= 16'h0528;    16'd56447: out <= 16'h041E;
    16'd56448: out <= 16'h0456;    16'd56449: out <= 16'hFE54;    16'd56450: out <= 16'h0180;    16'd56451: out <= 16'h013B;
    16'd56452: out <= 16'h0633;    16'd56453: out <= 16'h05C3;    16'd56454: out <= 16'h0814;    16'd56455: out <= 16'h0518;
    16'd56456: out <= 16'h0C01;    16'd56457: out <= 16'h00E3;    16'd56458: out <= 16'h05C0;    16'd56459: out <= 16'h0A53;
    16'd56460: out <= 16'h0631;    16'd56461: out <= 16'hFE8A;    16'd56462: out <= 16'hFF0D;    16'd56463: out <= 16'hFF72;
    16'd56464: out <= 16'h0077;    16'd56465: out <= 16'h06DD;    16'd56466: out <= 16'h0316;    16'd56467: out <= 16'h04F7;
    16'd56468: out <= 16'h009F;    16'd56469: out <= 16'h04DB;    16'd56470: out <= 16'h0334;    16'd56471: out <= 16'h0401;
    16'd56472: out <= 16'h04D8;    16'd56473: out <= 16'hFEAA;    16'd56474: out <= 16'h01A1;    16'd56475: out <= 16'h07B5;
    16'd56476: out <= 16'h02BA;    16'd56477: out <= 16'h0000;    16'd56478: out <= 16'h0584;    16'd56479: out <= 16'h0420;
    16'd56480: out <= 16'h01F7;    16'd56481: out <= 16'h05B8;    16'd56482: out <= 16'hFD6B;    16'd56483: out <= 16'h03F1;
    16'd56484: out <= 16'h0741;    16'd56485: out <= 16'h0963;    16'd56486: out <= 16'h07F7;    16'd56487: out <= 16'h06AD;
    16'd56488: out <= 16'hFD7F;    16'd56489: out <= 16'h0578;    16'd56490: out <= 16'hFF4C;    16'd56491: out <= 16'hFF63;
    16'd56492: out <= 16'h09BE;    16'd56493: out <= 16'h082A;    16'd56494: out <= 16'hFB5E;    16'd56495: out <= 16'hFEE7;
    16'd56496: out <= 16'h0293;    16'd56497: out <= 16'hFF20;    16'd56498: out <= 16'h0058;    16'd56499: out <= 16'h0794;
    16'd56500: out <= 16'h07EB;    16'd56501: out <= 16'h0252;    16'd56502: out <= 16'h0C2D;    16'd56503: out <= 16'h05FD;
    16'd56504: out <= 16'hFF97;    16'd56505: out <= 16'h06C4;    16'd56506: out <= 16'h0494;    16'd56507: out <= 16'hFB6B;
    16'd56508: out <= 16'h08BC;    16'd56509: out <= 16'h0288;    16'd56510: out <= 16'h04D0;    16'd56511: out <= 16'h074D;
    16'd56512: out <= 16'hFC09;    16'd56513: out <= 16'h01A2;    16'd56514: out <= 16'hFFE4;    16'd56515: out <= 16'h01B2;
    16'd56516: out <= 16'h0179;    16'd56517: out <= 16'hFA9A;    16'd56518: out <= 16'h028A;    16'd56519: out <= 16'h016F;
    16'd56520: out <= 16'h03D9;    16'd56521: out <= 16'h04E0;    16'd56522: out <= 16'h0067;    16'd56523: out <= 16'hFD61;
    16'd56524: out <= 16'h0F12;    16'd56525: out <= 16'h0108;    16'd56526: out <= 16'hFBF6;    16'd56527: out <= 16'hFE3B;
    16'd56528: out <= 16'hFEBD;    16'd56529: out <= 16'hFEF4;    16'd56530: out <= 16'h0449;    16'd56531: out <= 16'h01AB;
    16'd56532: out <= 16'hFE84;    16'd56533: out <= 16'h03A2;    16'd56534: out <= 16'hFE2C;    16'd56535: out <= 16'h0162;
    16'd56536: out <= 16'h0557;    16'd56537: out <= 16'hFDC3;    16'd56538: out <= 16'h0153;    16'd56539: out <= 16'hFF7C;
    16'd56540: out <= 16'h0006;    16'd56541: out <= 16'hFFEA;    16'd56542: out <= 16'hFD61;    16'd56543: out <= 16'hF9D0;
    16'd56544: out <= 16'hFF12;    16'd56545: out <= 16'hFC62;    16'd56546: out <= 16'hFF15;    16'd56547: out <= 16'h009E;
    16'd56548: out <= 16'hFD89;    16'd56549: out <= 16'hF9C2;    16'd56550: out <= 16'h04D1;    16'd56551: out <= 16'h042F;
    16'd56552: out <= 16'hFE1D;    16'd56553: out <= 16'h02D9;    16'd56554: out <= 16'hFB22;    16'd56555: out <= 16'h06B0;
    16'd56556: out <= 16'hFE29;    16'd56557: out <= 16'hFC19;    16'd56558: out <= 16'h0528;    16'd56559: out <= 16'h0203;
    16'd56560: out <= 16'hFB6F;    16'd56561: out <= 16'hFA11;    16'd56562: out <= 16'hFC60;    16'd56563: out <= 16'h0474;
    16'd56564: out <= 16'hFDC3;    16'd56565: out <= 16'hFD08;    16'd56566: out <= 16'h00EA;    16'd56567: out <= 16'hFA1F;
    16'd56568: out <= 16'hFBF1;    16'd56569: out <= 16'hFD50;    16'd56570: out <= 16'hFCE1;    16'd56571: out <= 16'h02A4;
    16'd56572: out <= 16'h0279;    16'd56573: out <= 16'h0046;    16'd56574: out <= 16'h0408;    16'd56575: out <= 16'hF8B6;
    16'd56576: out <= 16'h0452;    16'd56577: out <= 16'hFDBE;    16'd56578: out <= 16'h0859;    16'd56579: out <= 16'hFB9E;
    16'd56580: out <= 16'hFD11;    16'd56581: out <= 16'hFC17;    16'd56582: out <= 16'h0241;    16'd56583: out <= 16'hFFC4;
    16'd56584: out <= 16'h027C;    16'd56585: out <= 16'hFCDC;    16'd56586: out <= 16'hFE69;    16'd56587: out <= 16'hFB39;
    16'd56588: out <= 16'hFE1E;    16'd56589: out <= 16'h0739;    16'd56590: out <= 16'hF891;    16'd56591: out <= 16'h0482;
    16'd56592: out <= 16'h0316;    16'd56593: out <= 16'hFA46;    16'd56594: out <= 16'hF8D4;    16'd56595: out <= 16'h087A;
    16'd56596: out <= 16'h033F;    16'd56597: out <= 16'hFE59;    16'd56598: out <= 16'h02A0;    16'd56599: out <= 16'h024B;
    16'd56600: out <= 16'h050A;    16'd56601: out <= 16'hF803;    16'd56602: out <= 16'h03FB;    16'd56603: out <= 16'h07D6;
    16'd56604: out <= 16'h0207;    16'd56605: out <= 16'hFC65;    16'd56606: out <= 16'hFF46;    16'd56607: out <= 16'h014F;
    16'd56608: out <= 16'hFD53;    16'd56609: out <= 16'hF904;    16'd56610: out <= 16'hFCCF;    16'd56611: out <= 16'hFBB7;
    16'd56612: out <= 16'h00D2;    16'd56613: out <= 16'h0032;    16'd56614: out <= 16'h016A;    16'd56615: out <= 16'hF8D6;
    16'd56616: out <= 16'h00D7;    16'd56617: out <= 16'hFF1B;    16'd56618: out <= 16'hFE09;    16'd56619: out <= 16'h0142;
    16'd56620: out <= 16'hF773;    16'd56621: out <= 16'hFFFD;    16'd56622: out <= 16'hF709;    16'd56623: out <= 16'hFB12;
    16'd56624: out <= 16'h01DB;    16'd56625: out <= 16'h0B37;    16'd56626: out <= 16'h0993;    16'd56627: out <= 16'h0379;
    16'd56628: out <= 16'h078F;    16'd56629: out <= 16'hFCDD;    16'd56630: out <= 16'h0145;    16'd56631: out <= 16'hFF36;
    16'd56632: out <= 16'hFFC4;    16'd56633: out <= 16'h08B6;    16'd56634: out <= 16'h09A9;    16'd56635: out <= 16'h04F6;
    16'd56636: out <= 16'h01D0;    16'd56637: out <= 16'h06A2;    16'd56638: out <= 16'h000A;    16'd56639: out <= 16'h08EE;
    16'd56640: out <= 16'h025B;    16'd56641: out <= 16'h0458;    16'd56642: out <= 16'h0671;    16'd56643: out <= 16'h03B9;
    16'd56644: out <= 16'h05EB;    16'd56645: out <= 16'h00ED;    16'd56646: out <= 16'h0678;    16'd56647: out <= 16'h030A;
    16'd56648: out <= 16'h066A;    16'd56649: out <= 16'h0127;    16'd56650: out <= 16'hFEA8;    16'd56651: out <= 16'h059A;
    16'd56652: out <= 16'h040D;    16'd56653: out <= 16'h06D9;    16'd56654: out <= 16'h047A;    16'd56655: out <= 16'h074E;
    16'd56656: out <= 16'h0738;    16'd56657: out <= 16'h0339;    16'd56658: out <= 16'h02AD;    16'd56659: out <= 16'h015B;
    16'd56660: out <= 16'h0583;    16'd56661: out <= 16'h07D2;    16'd56662: out <= 16'hFF20;    16'd56663: out <= 16'h0BC3;
    16'd56664: out <= 16'h0490;    16'd56665: out <= 16'h034C;    16'd56666: out <= 16'hFBB6;    16'd56667: out <= 16'h09A5;
    16'd56668: out <= 16'h0297;    16'd56669: out <= 16'hFF86;    16'd56670: out <= 16'h027B;    16'd56671: out <= 16'h040C;
    16'd56672: out <= 16'hFC49;    16'd56673: out <= 16'h0790;    16'd56674: out <= 16'h06E2;    16'd56675: out <= 16'h0681;
    16'd56676: out <= 16'h06BD;    16'd56677: out <= 16'h081D;    16'd56678: out <= 16'h077F;    16'd56679: out <= 16'h07AC;
    16'd56680: out <= 16'h049C;    16'd56681: out <= 16'h012F;    16'd56682: out <= 16'h0628;    16'd56683: out <= 16'h0A26;
    16'd56684: out <= 16'hFF46;    16'd56685: out <= 16'h028B;    16'd56686: out <= 16'h0053;    16'd56687: out <= 16'h036C;
    16'd56688: out <= 16'h02DF;    16'd56689: out <= 16'hFEC4;    16'd56690: out <= 16'h0722;    16'd56691: out <= 16'h04B1;
    16'd56692: out <= 16'h0324;    16'd56693: out <= 16'h0884;    16'd56694: out <= 16'hFD98;    16'd56695: out <= 16'h0494;
    16'd56696: out <= 16'hFC07;    16'd56697: out <= 16'h07F9;    16'd56698: out <= 16'h0416;    16'd56699: out <= 16'h0829;
    16'd56700: out <= 16'h02CA;    16'd56701: out <= 16'h00BB;    16'd56702: out <= 16'h00FF;    16'd56703: out <= 16'h071E;
    16'd56704: out <= 16'h04B6;    16'd56705: out <= 16'h009D;    16'd56706: out <= 16'h073C;    16'd56707: out <= 16'h01BA;
    16'd56708: out <= 16'h0811;    16'd56709: out <= 16'h03C7;    16'd56710: out <= 16'h0014;    16'd56711: out <= 16'h0694;
    16'd56712: out <= 16'h0009;    16'd56713: out <= 16'h04D8;    16'd56714: out <= 16'hFF70;    16'd56715: out <= 16'h0399;
    16'd56716: out <= 16'hFE64;    16'd56717: out <= 16'h05A9;    16'd56718: out <= 16'h026A;    16'd56719: out <= 16'hFE1E;
    16'd56720: out <= 16'hFDB8;    16'd56721: out <= 16'hFFB6;    16'd56722: out <= 16'hFF90;    16'd56723: out <= 16'hFE78;
    16'd56724: out <= 16'hFBD9;    16'd56725: out <= 16'h0364;    16'd56726: out <= 16'hFE9E;    16'd56727: out <= 16'h063F;
    16'd56728: out <= 16'h09AC;    16'd56729: out <= 16'h065D;    16'd56730: out <= 16'h09AF;    16'd56731: out <= 16'h0805;
    16'd56732: out <= 16'h08CE;    16'd56733: out <= 16'h001B;    16'd56734: out <= 16'h02DB;    16'd56735: out <= 16'h02F8;
    16'd56736: out <= 16'hFFB5;    16'd56737: out <= 16'h0ABE;    16'd56738: out <= 16'hFE44;    16'd56739: out <= 16'h018F;
    16'd56740: out <= 16'h038B;    16'd56741: out <= 16'h0848;    16'd56742: out <= 16'h0CE6;    16'd56743: out <= 16'h0954;
    16'd56744: out <= 16'h0218;    16'd56745: out <= 16'h05BF;    16'd56746: out <= 16'h070C;    16'd56747: out <= 16'hFEA2;
    16'd56748: out <= 16'h0375;    16'd56749: out <= 16'h04B8;    16'd56750: out <= 16'h0169;    16'd56751: out <= 16'h0519;
    16'd56752: out <= 16'hFC9A;    16'd56753: out <= 16'h076A;    16'd56754: out <= 16'h04DB;    16'd56755: out <= 16'hFFAB;
    16'd56756: out <= 16'h0224;    16'd56757: out <= 16'h01FA;    16'd56758: out <= 16'h03EC;    16'd56759: out <= 16'h04E3;
    16'd56760: out <= 16'hFA88;    16'd56761: out <= 16'h0399;    16'd56762: out <= 16'h06C6;    16'd56763: out <= 16'h0748;
    16'd56764: out <= 16'h09F2;    16'd56765: out <= 16'hFEF9;    16'd56766: out <= 16'h0256;    16'd56767: out <= 16'h001F;
    16'd56768: out <= 16'h056F;    16'd56769: out <= 16'h0B97;    16'd56770: out <= 16'h05E0;    16'd56771: out <= 16'h017B;
    16'd56772: out <= 16'h03FC;    16'd56773: out <= 16'hFE70;    16'd56774: out <= 16'h0350;    16'd56775: out <= 16'h041B;
    16'd56776: out <= 16'h03E9;    16'd56777: out <= 16'hFFEE;    16'd56778: out <= 16'hFF66;    16'd56779: out <= 16'hFD7E;
    16'd56780: out <= 16'h0960;    16'd56781: out <= 16'h0226;    16'd56782: out <= 16'hFDFC;    16'd56783: out <= 16'h08E7;
    16'd56784: out <= 16'hFE58;    16'd56785: out <= 16'hFE3E;    16'd56786: out <= 16'h0058;    16'd56787: out <= 16'h01A5;
    16'd56788: out <= 16'h012C;    16'd56789: out <= 16'h0314;    16'd56790: out <= 16'hFC7F;    16'd56791: out <= 16'hFB1B;
    16'd56792: out <= 16'h01AF;    16'd56793: out <= 16'hFC8C;    16'd56794: out <= 16'hF997;    16'd56795: out <= 16'h03D7;
    16'd56796: out <= 16'h0003;    16'd56797: out <= 16'hFFC4;    16'd56798: out <= 16'hFBEC;    16'd56799: out <= 16'h035F;
    16'd56800: out <= 16'h0494;    16'd56801: out <= 16'h01EE;    16'd56802: out <= 16'h023C;    16'd56803: out <= 16'hFD95;
    16'd56804: out <= 16'h0671;    16'd56805: out <= 16'h0286;    16'd56806: out <= 16'h0092;    16'd56807: out <= 16'h02F7;
    16'd56808: out <= 16'h01D9;    16'd56809: out <= 16'h0819;    16'd56810: out <= 16'h00E9;    16'd56811: out <= 16'hFCD8;
    16'd56812: out <= 16'h043E;    16'd56813: out <= 16'hFBFC;    16'd56814: out <= 16'hFC59;    16'd56815: out <= 16'h0052;
    16'd56816: out <= 16'hFD5A;    16'd56817: out <= 16'hF9A8;    16'd56818: out <= 16'h0159;    16'd56819: out <= 16'hFBA6;
    16'd56820: out <= 16'hFB5D;    16'd56821: out <= 16'hF7D6;    16'd56822: out <= 16'hFF67;    16'd56823: out <= 16'h033B;
    16'd56824: out <= 16'hFB3F;    16'd56825: out <= 16'hFB7D;    16'd56826: out <= 16'hFFBC;    16'd56827: out <= 16'h05DD;
    16'd56828: out <= 16'h047C;    16'd56829: out <= 16'hFFD3;    16'd56830: out <= 16'hFC98;    16'd56831: out <= 16'hFFCD;
    16'd56832: out <= 16'h0253;    16'd56833: out <= 16'h01EB;    16'd56834: out <= 16'h0024;    16'd56835: out <= 16'h0001;
    16'd56836: out <= 16'h0268;    16'd56837: out <= 16'hF8C5;    16'd56838: out <= 16'hF9A8;    16'd56839: out <= 16'h05C8;
    16'd56840: out <= 16'hFCEF;    16'd56841: out <= 16'h02FC;    16'd56842: out <= 16'hFCF1;    16'd56843: out <= 16'h0215;
    16'd56844: out <= 16'hFBDC;    16'd56845: out <= 16'hFCD8;    16'd56846: out <= 16'h02CE;    16'd56847: out <= 16'hFEFA;
    16'd56848: out <= 16'h04B5;    16'd56849: out <= 16'h078A;    16'd56850: out <= 16'hFF57;    16'd56851: out <= 16'h013A;
    16'd56852: out <= 16'h06C6;    16'd56853: out <= 16'hFEE6;    16'd56854: out <= 16'hFA53;    16'd56855: out <= 16'hFE25;
    16'd56856: out <= 16'h0215;    16'd56857: out <= 16'h0A9D;    16'd56858: out <= 16'h00A6;    16'd56859: out <= 16'hFD6A;
    16'd56860: out <= 16'h0368;    16'd56861: out <= 16'hFE3E;    16'd56862: out <= 16'h02CA;    16'd56863: out <= 16'h00A1;
    16'd56864: out <= 16'h00EA;    16'd56865: out <= 16'h0225;    16'd56866: out <= 16'hFFBE;    16'd56867: out <= 16'hF6FB;
    16'd56868: out <= 16'h01AB;    16'd56869: out <= 16'h01F3;    16'd56870: out <= 16'h0210;    16'd56871: out <= 16'h030B;
    16'd56872: out <= 16'hF8F0;    16'd56873: out <= 16'hFF9D;    16'd56874: out <= 16'h0099;    16'd56875: out <= 16'hFE55;
    16'd56876: out <= 16'h03A6;    16'd56877: out <= 16'hFB86;    16'd56878: out <= 16'h0144;    16'd56879: out <= 16'h0277;
    16'd56880: out <= 16'h03D0;    16'd56881: out <= 16'h09C4;    16'd56882: out <= 16'h0586;    16'd56883: out <= 16'h047A;
    16'd56884: out <= 16'h03D7;    16'd56885: out <= 16'h0329;    16'd56886: out <= 16'h0962;    16'd56887: out <= 16'h046E;
    16'd56888: out <= 16'h02D4;    16'd56889: out <= 16'h067A;    16'd56890: out <= 16'h05B6;    16'd56891: out <= 16'h006F;
    16'd56892: out <= 16'h01FF;    16'd56893: out <= 16'hFE6C;    16'd56894: out <= 16'hFCB3;    16'd56895: out <= 16'hFE82;
    16'd56896: out <= 16'h004D;    16'd56897: out <= 16'hFFF4;    16'd56898: out <= 16'h04E6;    16'd56899: out <= 16'h0414;
    16'd56900: out <= 16'h03AD;    16'd56901: out <= 16'h027A;    16'd56902: out <= 16'h07F1;    16'd56903: out <= 16'h0286;
    16'd56904: out <= 16'h02C9;    16'd56905: out <= 16'h008D;    16'd56906: out <= 16'h0284;    16'd56907: out <= 16'h0456;
    16'd56908: out <= 16'h046F;    16'd56909: out <= 16'h00A4;    16'd56910: out <= 16'h024E;    16'd56911: out <= 16'h01EC;
    16'd56912: out <= 16'h010F;    16'd56913: out <= 16'h012D;    16'd56914: out <= 16'h020B;    16'd56915: out <= 16'hFD6F;
    16'd56916: out <= 16'h05FD;    16'd56917: out <= 16'h0245;    16'd56918: out <= 16'hFB11;    16'd56919: out <= 16'h0404;
    16'd56920: out <= 16'h0755;    16'd56921: out <= 16'h0627;    16'd56922: out <= 16'h01CB;    16'd56923: out <= 16'hFEFC;
    16'd56924: out <= 16'h081F;    16'd56925: out <= 16'h0317;    16'd56926: out <= 16'h03E2;    16'd56927: out <= 16'h05E8;
    16'd56928: out <= 16'h030B;    16'd56929: out <= 16'h00F0;    16'd56930: out <= 16'h005D;    16'd56931: out <= 16'h083F;
    16'd56932: out <= 16'h084E;    16'd56933: out <= 16'hFE5A;    16'd56934: out <= 16'hFFD9;    16'd56935: out <= 16'h0302;
    16'd56936: out <= 16'h05B0;    16'd56937: out <= 16'h07C3;    16'd56938: out <= 16'hFFD9;    16'd56939: out <= 16'h0F17;
    16'd56940: out <= 16'h0203;    16'd56941: out <= 16'h02DD;    16'd56942: out <= 16'h009A;    16'd56943: out <= 16'h083D;
    16'd56944: out <= 16'h06CD;    16'd56945: out <= 16'h0414;    16'd56946: out <= 16'h0542;    16'd56947: out <= 16'h0180;
    16'd56948: out <= 16'h067D;    16'd56949: out <= 16'h029E;    16'd56950: out <= 16'h0028;    16'd56951: out <= 16'hFC65;
    16'd56952: out <= 16'h030A;    16'd56953: out <= 16'h0546;    16'd56954: out <= 16'h074C;    16'd56955: out <= 16'h0337;
    16'd56956: out <= 16'h059F;    16'd56957: out <= 16'h05F1;    16'd56958: out <= 16'h0688;    16'd56959: out <= 16'h01A8;
    16'd56960: out <= 16'h0176;    16'd56961: out <= 16'h00A0;    16'd56962: out <= 16'hFF09;    16'd56963: out <= 16'h0650;
    16'd56964: out <= 16'h0631;    16'd56965: out <= 16'h0644;    16'd56966: out <= 16'h088A;    16'd56967: out <= 16'h0298;
    16'd56968: out <= 16'h0621;    16'd56969: out <= 16'h03D4;    16'd56970: out <= 16'h03B4;    16'd56971: out <= 16'h05F1;
    16'd56972: out <= 16'hFE1C;    16'd56973: out <= 16'h0582;    16'd56974: out <= 16'hFEA1;    16'd56975: out <= 16'h04D4;
    16'd56976: out <= 16'h0848;    16'd56977: out <= 16'h0B4B;    16'd56978: out <= 16'h007D;    16'd56979: out <= 16'h09E9;
    16'd56980: out <= 16'h00C3;    16'd56981: out <= 16'h06A4;    16'd56982: out <= 16'h0231;    16'd56983: out <= 16'h07BA;
    16'd56984: out <= 16'hFFC7;    16'd56985: out <= 16'h01F3;    16'd56986: out <= 16'h024A;    16'd56987: out <= 16'h025A;
    16'd56988: out <= 16'h0440;    16'd56989: out <= 16'h0892;    16'd56990: out <= 16'hFEB1;    16'd56991: out <= 16'hFCD7;
    16'd56992: out <= 16'h05E3;    16'd56993: out <= 16'h0538;    16'd56994: out <= 16'h028B;    16'd56995: out <= 16'h010F;
    16'd56996: out <= 16'h0715;    16'd56997: out <= 16'h0581;    16'd56998: out <= 16'h07CB;    16'd56999: out <= 16'h0585;
    16'd57000: out <= 16'h0611;    16'd57001: out <= 16'h0873;    16'd57002: out <= 16'h0325;    16'd57003: out <= 16'hFE76;
    16'd57004: out <= 16'hFFC7;    16'd57005: out <= 16'h0636;    16'd57006: out <= 16'hFFF6;    16'd57007: out <= 16'h00ED;
    16'd57008: out <= 16'h0170;    16'd57009: out <= 16'h01FB;    16'd57010: out <= 16'h0434;    16'd57011: out <= 16'h0752;
    16'd57012: out <= 16'h03DF;    16'd57013: out <= 16'h0570;    16'd57014: out <= 16'hFDDC;    16'd57015: out <= 16'h020F;
    16'd57016: out <= 16'h07EA;    16'd57017: out <= 16'h026B;    16'd57018: out <= 16'h0AC5;    16'd57019: out <= 16'h0614;
    16'd57020: out <= 16'hFF5D;    16'd57021: out <= 16'h03E3;    16'd57022: out <= 16'h0444;    16'd57023: out <= 16'h0413;
    16'd57024: out <= 16'h0713;    16'd57025: out <= 16'h0538;    16'd57026: out <= 16'hFEC8;    16'd57027: out <= 16'hFF62;
    16'd57028: out <= 16'hFE70;    16'd57029: out <= 16'hFEBC;    16'd57030: out <= 16'h01C1;    16'd57031: out <= 16'h0275;
    16'd57032: out <= 16'hFE34;    16'd57033: out <= 16'hFE34;    16'd57034: out <= 16'hFA11;    16'd57035: out <= 16'h0076;
    16'd57036: out <= 16'hFB3E;    16'd57037: out <= 16'h0332;    16'd57038: out <= 16'hFFBF;    16'd57039: out <= 16'hFDA1;
    16'd57040: out <= 16'h0608;    16'd57041: out <= 16'h002A;    16'd57042: out <= 16'h012D;    16'd57043: out <= 16'hFF72;
    16'd57044: out <= 16'hFDD6;    16'd57045: out <= 16'hFD66;    16'd57046: out <= 16'hF7B3;    16'd57047: out <= 16'h081A;
    16'd57048: out <= 16'h05EB;    16'd57049: out <= 16'hF90B;    16'd57050: out <= 16'hFEE7;    16'd57051: out <= 16'h03E8;
    16'd57052: out <= 16'hFE09;    16'd57053: out <= 16'h0443;    16'd57054: out <= 16'hFC6C;    16'd57055: out <= 16'hFA6E;
    16'd57056: out <= 16'hFE1A;    16'd57057: out <= 16'h05FD;    16'd57058: out <= 16'h0517;    16'd57059: out <= 16'hFFAC;
    16'd57060: out <= 16'h02CE;    16'd57061: out <= 16'h01F0;    16'd57062: out <= 16'hFF17;    16'd57063: out <= 16'hFD68;
    16'd57064: out <= 16'h004E;    16'd57065: out <= 16'hFD87;    16'd57066: out <= 16'hFC1D;    16'd57067: out <= 16'h0352;
    16'd57068: out <= 16'h0134;    16'd57069: out <= 16'h0120;    16'd57070: out <= 16'hFD3E;    16'd57071: out <= 16'h03D5;
    16'd57072: out <= 16'h0018;    16'd57073: out <= 16'h0076;    16'd57074: out <= 16'h02C2;    16'd57075: out <= 16'hFDC3;
    16'd57076: out <= 16'h02AB;    16'd57077: out <= 16'h044E;    16'd57078: out <= 16'hFDF6;    16'd57079: out <= 16'hFF8A;
    16'd57080: out <= 16'h04AE;    16'd57081: out <= 16'h0118;    16'd57082: out <= 16'hFD9C;    16'd57083: out <= 16'hFF8D;
    16'd57084: out <= 16'h01E2;    16'd57085: out <= 16'hFFDD;    16'd57086: out <= 16'h00F2;    16'd57087: out <= 16'h0673;
    16'd57088: out <= 16'h01E1;    16'd57089: out <= 16'h006F;    16'd57090: out <= 16'h06D9;    16'd57091: out <= 16'hFDC2;
    16'd57092: out <= 16'hFE10;    16'd57093: out <= 16'h05AD;    16'd57094: out <= 16'h017D;    16'd57095: out <= 16'h01D0;
    16'd57096: out <= 16'h04E8;    16'd57097: out <= 16'hFD5A;    16'd57098: out <= 16'hFEF1;    16'd57099: out <= 16'hFE87;
    16'd57100: out <= 16'h04D7;    16'd57101: out <= 16'hFD31;    16'd57102: out <= 16'hFF5F;    16'd57103: out <= 16'hFCDC;
    16'd57104: out <= 16'h024E;    16'd57105: out <= 16'h0305;    16'd57106: out <= 16'h0376;    16'd57107: out <= 16'h06FD;
    16'd57108: out <= 16'hF686;    16'd57109: out <= 16'hFB4F;    16'd57110: out <= 16'hFF13;    16'd57111: out <= 16'hFA68;
    16'd57112: out <= 16'h07AB;    16'd57113: out <= 16'hFDB0;    16'd57114: out <= 16'hFA61;    16'd57115: out <= 16'hF75E;
    16'd57116: out <= 16'h029E;    16'd57117: out <= 16'hFE80;    16'd57118: out <= 16'h00EE;    16'd57119: out <= 16'h0427;
    16'd57120: out <= 16'h003A;    16'd57121: out <= 16'hFDFD;    16'd57122: out <= 16'h00FD;    16'd57123: out <= 16'h0161;
    16'd57124: out <= 16'h04AB;    16'd57125: out <= 16'hF9A3;    16'd57126: out <= 16'h0501;    16'd57127: out <= 16'h0003;
    16'd57128: out <= 16'hFF0B;    16'd57129: out <= 16'hFB04;    16'd57130: out <= 16'h002E;    16'd57131: out <= 16'hF4F6;
    16'd57132: out <= 16'hF98C;    16'd57133: out <= 16'h03B3;    16'd57134: out <= 16'h0007;    16'd57135: out <= 16'hF943;
    16'd57136: out <= 16'hFCF8;    16'd57137: out <= 16'h0BE2;    16'd57138: out <= 16'h011C;    16'd57139: out <= 16'h03AC;
    16'd57140: out <= 16'h0055;    16'd57141: out <= 16'h0080;    16'd57142: out <= 16'h00AC;    16'd57143: out <= 16'h03B5;
    16'd57144: out <= 16'h0607;    16'd57145: out <= 16'h03EC;    16'd57146: out <= 16'h03E9;    16'd57147: out <= 16'h086E;
    16'd57148: out <= 16'h0029;    16'd57149: out <= 16'h023B;    16'd57150: out <= 16'h031E;    16'd57151: out <= 16'h05D5;
    16'd57152: out <= 16'h0BFE;    16'd57153: out <= 16'h02DC;    16'd57154: out <= 16'h065D;    16'd57155: out <= 16'hFE11;
    16'd57156: out <= 16'h0583;    16'd57157: out <= 16'h0C6B;    16'd57158: out <= 16'h0095;    16'd57159: out <= 16'h02D3;
    16'd57160: out <= 16'h0549;    16'd57161: out <= 16'h0338;    16'd57162: out <= 16'h0343;    16'd57163: out <= 16'hFE15;
    16'd57164: out <= 16'h04EB;    16'd57165: out <= 16'h0547;    16'd57166: out <= 16'h0645;    16'd57167: out <= 16'h05A4;
    16'd57168: out <= 16'h0672;    16'd57169: out <= 16'h00B7;    16'd57170: out <= 16'hFF29;    16'd57171: out <= 16'h0AA8;
    16'd57172: out <= 16'h0381;    16'd57173: out <= 16'h059E;    16'd57174: out <= 16'h041D;    16'd57175: out <= 16'hFEC2;
    16'd57176: out <= 16'h04E1;    16'd57177: out <= 16'h024B;    16'd57178: out <= 16'h02FD;    16'd57179: out <= 16'h0C0A;
    16'd57180: out <= 16'h0B0E;    16'd57181: out <= 16'h0027;    16'd57182: out <= 16'h076E;    16'd57183: out <= 16'h059E;
    16'd57184: out <= 16'h05CD;    16'd57185: out <= 16'h017A;    16'd57186: out <= 16'h07D7;    16'd57187: out <= 16'h0350;
    16'd57188: out <= 16'h00DE;    16'd57189: out <= 16'h03A3;    16'd57190: out <= 16'h00FF;    16'd57191: out <= 16'h06C1;
    16'd57192: out <= 16'h0ACF;    16'd57193: out <= 16'h09C2;    16'd57194: out <= 16'hFC1E;    16'd57195: out <= 16'h0947;
    16'd57196: out <= 16'h04D7;    16'd57197: out <= 16'h04EC;    16'd57198: out <= 16'h013D;    16'd57199: out <= 16'h0620;
    16'd57200: out <= 16'h0A09;    16'd57201: out <= 16'h00E4;    16'd57202: out <= 16'h03CE;    16'd57203: out <= 16'h0219;
    16'd57204: out <= 16'h0C16;    16'd57205: out <= 16'h0259;    16'd57206: out <= 16'hFDF0;    16'd57207: out <= 16'h04C6;
    16'd57208: out <= 16'h08B6;    16'd57209: out <= 16'h01FB;    16'd57210: out <= 16'h05B2;    16'd57211: out <= 16'h0703;
    16'd57212: out <= 16'h0921;    16'd57213: out <= 16'hFF2D;    16'd57214: out <= 16'h0C36;    16'd57215: out <= 16'h0713;
    16'd57216: out <= 16'h0318;    16'd57217: out <= 16'hFD91;    16'd57218: out <= 16'h07B4;    16'd57219: out <= 16'hFCE5;
    16'd57220: out <= 16'h0923;    16'd57221: out <= 16'h092E;    16'd57222: out <= 16'h012C;    16'd57223: out <= 16'h038E;
    16'd57224: out <= 16'h022D;    16'd57225: out <= 16'h0730;    16'd57226: out <= 16'h07D5;    16'd57227: out <= 16'h04C9;
    16'd57228: out <= 16'h0C79;    16'd57229: out <= 16'h00B2;    16'd57230: out <= 16'h0744;    16'd57231: out <= 16'h04EE;
    16'd57232: out <= 16'h06B7;    16'd57233: out <= 16'hFD5D;    16'd57234: out <= 16'h0267;    16'd57235: out <= 16'h02F2;
    16'd57236: out <= 16'h01C7;    16'd57237: out <= 16'h002D;    16'd57238: out <= 16'h04DC;    16'd57239: out <= 16'h0566;
    16'd57240: out <= 16'h0364;    16'd57241: out <= 16'h05A1;    16'd57242: out <= 16'h023A;    16'd57243: out <= 16'h030D;
    16'd57244: out <= 16'h053C;    16'd57245: out <= 16'h007B;    16'd57246: out <= 16'h068F;    16'd57247: out <= 16'h02F8;
    16'd57248: out <= 16'h0653;    16'd57249: out <= 16'h0B19;    16'd57250: out <= 16'h0A00;    16'd57251: out <= 16'h0604;
    16'd57252: out <= 16'h066F;    16'd57253: out <= 16'h02C4;    16'd57254: out <= 16'h0E46;    16'd57255: out <= 16'h0944;
    16'd57256: out <= 16'h056F;    16'd57257: out <= 16'h0384;    16'd57258: out <= 16'hFF2E;    16'd57259: out <= 16'h01FB;
    16'd57260: out <= 16'h0205;    16'd57261: out <= 16'h06BB;    16'd57262: out <= 16'h050E;    16'd57263: out <= 16'h03A2;
    16'd57264: out <= 16'h04DC;    16'd57265: out <= 16'h0513;    16'd57266: out <= 16'h0A94;    16'd57267: out <= 16'hFCCD;
    16'd57268: out <= 16'h0B9B;    16'd57269: out <= 16'h03CA;    16'd57270: out <= 16'h07F9;    16'd57271: out <= 16'hFF6E;
    16'd57272: out <= 16'hFE9B;    16'd57273: out <= 16'h001C;    16'd57274: out <= 16'h04DE;    16'd57275: out <= 16'h0443;
    16'd57276: out <= 16'h0601;    16'd57277: out <= 16'h033C;    16'd57278: out <= 16'h029A;    16'd57279: out <= 16'h01A2;
    16'd57280: out <= 16'h045C;    16'd57281: out <= 16'h0984;    16'd57282: out <= 16'h045A;    16'd57283: out <= 16'hFB50;
    16'd57284: out <= 16'h057A;    16'd57285: out <= 16'h00B9;    16'd57286: out <= 16'h028E;    16'd57287: out <= 16'hFC89;
    16'd57288: out <= 16'hF56F;    16'd57289: out <= 16'h03BE;    16'd57290: out <= 16'hF8BF;    16'd57291: out <= 16'h035F;
    16'd57292: out <= 16'hFEFA;    16'd57293: out <= 16'hFCA8;    16'd57294: out <= 16'h02E9;    16'd57295: out <= 16'hFBB8;
    16'd57296: out <= 16'h05CC;    16'd57297: out <= 16'h06BC;    16'd57298: out <= 16'hFD97;    16'd57299: out <= 16'hFBE6;
    16'd57300: out <= 16'h0094;    16'd57301: out <= 16'h0592;    16'd57302: out <= 16'h052D;    16'd57303: out <= 16'hFE11;
    16'd57304: out <= 16'h00DD;    16'd57305: out <= 16'h04B9;    16'd57306: out <= 16'hFF44;    16'd57307: out <= 16'hFEDC;
    16'd57308: out <= 16'h009B;    16'd57309: out <= 16'h0701;    16'd57310: out <= 16'hFA36;    16'd57311: out <= 16'hFF5B;
    16'd57312: out <= 16'hFAC1;    16'd57313: out <= 16'h02CA;    16'd57314: out <= 16'hFFCB;    16'd57315: out <= 16'hFF95;
    16'd57316: out <= 16'hFC4C;    16'd57317: out <= 16'hFBAE;    16'd57318: out <= 16'h07D3;    16'd57319: out <= 16'hF838;
    16'd57320: out <= 16'hFC3A;    16'd57321: out <= 16'h0304;    16'd57322: out <= 16'hFD7E;    16'd57323: out <= 16'h03C3;
    16'd57324: out <= 16'h03AD;    16'd57325: out <= 16'hFF77;    16'd57326: out <= 16'hFDEE;    16'd57327: out <= 16'hFAC7;
    16'd57328: out <= 16'h01EA;    16'd57329: out <= 16'hF94B;    16'd57330: out <= 16'hFB5C;    16'd57331: out <= 16'h02CE;
    16'd57332: out <= 16'h05A1;    16'd57333: out <= 16'hFF09;    16'd57334: out <= 16'h0249;    16'd57335: out <= 16'h0362;
    16'd57336: out <= 16'h01EF;    16'd57337: out <= 16'h00AE;    16'd57338: out <= 16'hFF68;    16'd57339: out <= 16'hFC07;
    16'd57340: out <= 16'h02BC;    16'd57341: out <= 16'hFECC;    16'd57342: out <= 16'hFC92;    16'd57343: out <= 16'h0499;
    16'd57344: out <= 16'hFBF5;    16'd57345: out <= 16'h062C;    16'd57346: out <= 16'h0256;    16'd57347: out <= 16'hF9F0;
    16'd57348: out <= 16'hF9ED;    16'd57349: out <= 16'h005F;    16'd57350: out <= 16'h01E6;    16'd57351: out <= 16'h0062;
    16'd57352: out <= 16'hFECC;    16'd57353: out <= 16'h0146;    16'd57354: out <= 16'h0597;    16'd57355: out <= 16'h03CC;
    16'd57356: out <= 16'h0163;    16'd57357: out <= 16'h022D;    16'd57358: out <= 16'h061B;    16'd57359: out <= 16'h02FC;
    16'd57360: out <= 16'hFAA0;    16'd57361: out <= 16'hFE96;    16'd57362: out <= 16'hFC84;    16'd57363: out <= 16'hF9E1;
    16'd57364: out <= 16'hF5CB;    16'd57365: out <= 16'hFD25;    16'd57366: out <= 16'hFCC0;    16'd57367: out <= 16'hF947;
    16'd57368: out <= 16'hFFC7;    16'd57369: out <= 16'h07CC;    16'd57370: out <= 16'h016B;    16'd57371: out <= 16'h01BC;
    16'd57372: out <= 16'h04E4;    16'd57373: out <= 16'hFB74;    16'd57374: out <= 16'h015E;    16'd57375: out <= 16'h0671;
    16'd57376: out <= 16'h00BA;    16'd57377: out <= 16'hFBA0;    16'd57378: out <= 16'hFF4A;    16'd57379: out <= 16'hFE0E;
    16'd57380: out <= 16'hFCA9;    16'd57381: out <= 16'h02AB;    16'd57382: out <= 16'hFCE9;    16'd57383: out <= 16'hFADF;
    16'd57384: out <= 16'h029D;    16'd57385: out <= 16'h00BA;    16'd57386: out <= 16'hFB43;    16'd57387: out <= 16'h010C;
    16'd57388: out <= 16'h0174;    16'd57389: out <= 16'h0078;    16'd57390: out <= 16'h0172;    16'd57391: out <= 16'h0236;
    16'd57392: out <= 16'h07BD;    16'd57393: out <= 16'h0578;    16'd57394: out <= 16'h081B;    16'd57395: out <= 16'h0219;
    16'd57396: out <= 16'hFECF;    16'd57397: out <= 16'h0257;    16'd57398: out <= 16'h0B23;    16'd57399: out <= 16'h0458;
    16'd57400: out <= 16'h0974;    16'd57401: out <= 16'h02D4;    16'd57402: out <= 16'hFDB6;    16'd57403: out <= 16'hF9AC;
    16'd57404: out <= 16'h02A2;    16'd57405: out <= 16'h06CE;    16'd57406: out <= 16'h041F;    16'd57407: out <= 16'h0836;
    16'd57408: out <= 16'h04C0;    16'd57409: out <= 16'h0743;    16'd57410: out <= 16'h0A90;    16'd57411: out <= 16'h0485;
    16'd57412: out <= 16'h0162;    16'd57413: out <= 16'h0186;    16'd57414: out <= 16'h0124;    16'd57415: out <= 16'hFFE4;
    16'd57416: out <= 16'h042D;    16'd57417: out <= 16'h0B5B;    16'd57418: out <= 16'h04C1;    16'd57419: out <= 16'hFF76;
    16'd57420: out <= 16'h0782;    16'd57421: out <= 16'h00FA;    16'd57422: out <= 16'h0764;    16'd57423: out <= 16'h02A8;
    16'd57424: out <= 16'h0403;    16'd57425: out <= 16'hFF27;    16'd57426: out <= 16'h05F8;    16'd57427: out <= 16'h0ABB;
    16'd57428: out <= 16'h010C;    16'd57429: out <= 16'h06C5;    16'd57430: out <= 16'h03CC;    16'd57431: out <= 16'h066B;
    16'd57432: out <= 16'h0259;    16'd57433: out <= 16'h0105;    16'd57434: out <= 16'hFF0F;    16'd57435: out <= 16'hFCAC;
    16'd57436: out <= 16'h06ED;    16'd57437: out <= 16'h02AE;    16'd57438: out <= 16'hFFA5;    16'd57439: out <= 16'hFCA3;
    16'd57440: out <= 16'h0132;    16'd57441: out <= 16'h0311;    16'd57442: out <= 16'h0F22;    16'd57443: out <= 16'h0863;
    16'd57444: out <= 16'h08E8;    16'd57445: out <= 16'hFEE7;    16'd57446: out <= 16'h0451;    16'd57447: out <= 16'h0A61;
    16'd57448: out <= 16'h049A;    16'd57449: out <= 16'h075E;    16'd57450: out <= 16'h0563;    16'd57451: out <= 16'h0337;
    16'd57452: out <= 16'h01EB;    16'd57453: out <= 16'h03F5;    16'd57454: out <= 16'h0A0D;    16'd57455: out <= 16'h09BC;
    16'd57456: out <= 16'h06C0;    16'd57457: out <= 16'h04BF;    16'd57458: out <= 16'h058E;    16'd57459: out <= 16'h07CC;
    16'd57460: out <= 16'h01DC;    16'd57461: out <= 16'h0126;    16'd57462: out <= 16'hFC1D;    16'd57463: out <= 16'h036F;
    16'd57464: out <= 16'hFFBD;    16'd57465: out <= 16'h062F;    16'd57466: out <= 16'h00E5;    16'd57467: out <= 16'h0803;
    16'd57468: out <= 16'h0776;    16'd57469: out <= 16'h01E1;    16'd57470: out <= 16'h0650;    16'd57471: out <= 16'h07FC;
    16'd57472: out <= 16'h01E0;    16'd57473: out <= 16'h0400;    16'd57474: out <= 16'h046A;    16'd57475: out <= 16'h0376;
    16'd57476: out <= 16'h002A;    16'd57477: out <= 16'h0860;    16'd57478: out <= 16'h045C;    16'd57479: out <= 16'h0404;
    16'd57480: out <= 16'h0BF9;    16'd57481: out <= 16'h023C;    16'd57482: out <= 16'h061F;    16'd57483: out <= 16'h019D;
    16'd57484: out <= 16'h0128;    16'd57485: out <= 16'h06DE;    16'd57486: out <= 16'h0387;    16'd57487: out <= 16'h00AD;
    16'd57488: out <= 16'h087E;    16'd57489: out <= 16'hFFAC;    16'd57490: out <= 16'hFC2D;    16'd57491: out <= 16'h0719;
    16'd57492: out <= 16'h08E1;    16'd57493: out <= 16'hFF64;    16'd57494: out <= 16'h06C0;    16'd57495: out <= 16'hF95D;
    16'd57496: out <= 16'h05A0;    16'd57497: out <= 16'h0458;    16'd57498: out <= 16'h04D4;    16'd57499: out <= 16'h0C01;
    16'd57500: out <= 16'h0378;    16'd57501: out <= 16'h07E8;    16'd57502: out <= 16'h097C;    16'd57503: out <= 16'h02BF;
    16'd57504: out <= 16'h00FC;    16'd57505: out <= 16'h056C;    16'd57506: out <= 16'h09FD;    16'd57507: out <= 16'h00AD;
    16'd57508: out <= 16'h011C;    16'd57509: out <= 16'h064B;    16'd57510: out <= 16'h05B3;    16'd57511: out <= 16'h0C30;
    16'd57512: out <= 16'h0A6D;    16'd57513: out <= 16'h0788;    16'd57514: out <= 16'h00DE;    16'd57515: out <= 16'hFFEF;
    16'd57516: out <= 16'h0740;    16'd57517: out <= 16'hFCC1;    16'd57518: out <= 16'h0144;    16'd57519: out <= 16'hFC89;
    16'd57520: out <= 16'h0535;    16'd57521: out <= 16'h0769;    16'd57522: out <= 16'hFE68;    16'd57523: out <= 16'h053A;
    16'd57524: out <= 16'h0733;    16'd57525: out <= 16'h0313;    16'd57526: out <= 16'h04F9;    16'd57527: out <= 16'h0547;
    16'd57528: out <= 16'h0B65;    16'd57529: out <= 16'h0978;    16'd57530: out <= 16'h0783;    16'd57531: out <= 16'h0084;
    16'd57532: out <= 16'h0AB4;    16'd57533: out <= 16'h04E3;    16'd57534: out <= 16'h055B;    16'd57535: out <= 16'h0158;
    16'd57536: out <= 16'h0A78;    16'd57537: out <= 16'h09A2;    16'd57538: out <= 16'hFA29;    16'd57539: out <= 16'h02C1;
    16'd57540: out <= 16'hFE43;    16'd57541: out <= 16'h031D;    16'd57542: out <= 16'hFF7B;    16'd57543: out <= 16'hFC69;
    16'd57544: out <= 16'hF9F9;    16'd57545: out <= 16'h0927;    16'd57546: out <= 16'hFF2E;    16'd57547: out <= 16'hFDDE;
    16'd57548: out <= 16'h0308;    16'd57549: out <= 16'h0D3E;    16'd57550: out <= 16'h02F1;    16'd57551: out <= 16'hFEA8;
    16'd57552: out <= 16'hFFD6;    16'd57553: out <= 16'hFEB9;    16'd57554: out <= 16'h07EA;    16'd57555: out <= 16'hF3B4;
    16'd57556: out <= 16'hF77B;    16'd57557: out <= 16'h04F1;    16'd57558: out <= 16'hFA8B;    16'd57559: out <= 16'h0583;
    16'd57560: out <= 16'hFF24;    16'd57561: out <= 16'hFAF9;    16'd57562: out <= 16'hFEC1;    16'd57563: out <= 16'hFF8D;
    16'd57564: out <= 16'hFFCC;    16'd57565: out <= 16'hFA4D;    16'd57566: out <= 16'hFAE9;    16'd57567: out <= 16'h0439;
    16'd57568: out <= 16'hFF54;    16'd57569: out <= 16'h03CC;    16'd57570: out <= 16'hFD75;    16'd57571: out <= 16'h065C;
    16'd57572: out <= 16'hFB11;    16'd57573: out <= 16'h0116;    16'd57574: out <= 16'h00DE;    16'd57575: out <= 16'h0168;
    16'd57576: out <= 16'h01B6;    16'd57577: out <= 16'hFEB0;    16'd57578: out <= 16'hFF53;    16'd57579: out <= 16'h052D;
    16'd57580: out <= 16'h0585;    16'd57581: out <= 16'hFB5D;    16'd57582: out <= 16'h00EA;    16'd57583: out <= 16'h0159;
    16'd57584: out <= 16'h0188;    16'd57585: out <= 16'hFF61;    16'd57586: out <= 16'h0276;    16'd57587: out <= 16'h01EC;
    16'd57588: out <= 16'hFE0A;    16'd57589: out <= 16'hFF7F;    16'd57590: out <= 16'hFAAE;    16'd57591: out <= 16'hFF43;
    16'd57592: out <= 16'hFD8E;    16'd57593: out <= 16'hFD10;    16'd57594: out <= 16'h07FF;    16'd57595: out <= 16'hF82F;
    16'd57596: out <= 16'h00D8;    16'd57597: out <= 16'hFF71;    16'd57598: out <= 16'h0249;    16'd57599: out <= 16'hFEFC;
    16'd57600: out <= 16'hFF0A;    16'd57601: out <= 16'hFD1F;    16'd57602: out <= 16'hFD54;    16'd57603: out <= 16'h0493;
    16'd57604: out <= 16'h0271;    16'd57605: out <= 16'hFEBB;    16'd57606: out <= 16'h02B4;    16'd57607: out <= 16'h0377;
    16'd57608: out <= 16'h0014;    16'd57609: out <= 16'hFB5A;    16'd57610: out <= 16'h0A57;    16'd57611: out <= 16'hFF31;
    16'd57612: out <= 16'h047F;    16'd57613: out <= 16'hF89F;    16'd57614: out <= 16'h049C;    16'd57615: out <= 16'hFFA5;
    16'd57616: out <= 16'hFCF2;    16'd57617: out <= 16'h0071;    16'd57618: out <= 16'h029C;    16'd57619: out <= 16'h01C1;
    16'd57620: out <= 16'hFE5B;    16'd57621: out <= 16'hFEC4;    16'd57622: out <= 16'hFDFB;    16'd57623: out <= 16'hF73F;
    16'd57624: out <= 16'h03A5;    16'd57625: out <= 16'hFEC9;    16'd57626: out <= 16'hFEBC;    16'd57627: out <= 16'h05F9;
    16'd57628: out <= 16'h03A4;    16'd57629: out <= 16'h05A6;    16'd57630: out <= 16'h02E5;    16'd57631: out <= 16'hFC42;
    16'd57632: out <= 16'hF996;    16'd57633: out <= 16'hFBFD;    16'd57634: out <= 16'h050B;    16'd57635: out <= 16'hF6B7;
    16'd57636: out <= 16'h01A0;    16'd57637: out <= 16'hFCF6;    16'd57638: out <= 16'h00B5;    16'd57639: out <= 16'hFDAE;
    16'd57640: out <= 16'hFFC0;    16'd57641: out <= 16'hFE48;    16'd57642: out <= 16'hFABF;    16'd57643: out <= 16'hFE11;
    16'd57644: out <= 16'h04B7;    16'd57645: out <= 16'h01BA;    16'd57646: out <= 16'hFEA4;    16'd57647: out <= 16'hFE29;
    16'd57648: out <= 16'h03F1;    16'd57649: out <= 16'h0548;    16'd57650: out <= 16'h05B4;    16'd57651: out <= 16'h088C;
    16'd57652: out <= 16'h03CB;    16'd57653: out <= 16'h07B4;    16'd57654: out <= 16'h0126;    16'd57655: out <= 16'h0732;
    16'd57656: out <= 16'h098B;    16'd57657: out <= 16'h0961;    16'd57658: out <= 16'h0954;    16'd57659: out <= 16'h0175;
    16'd57660: out <= 16'h00C7;    16'd57661: out <= 16'hFDFC;    16'd57662: out <= 16'h0661;    16'd57663: out <= 16'hFDCD;
    16'd57664: out <= 16'h030A;    16'd57665: out <= 16'h065D;    16'd57666: out <= 16'h0627;    16'd57667: out <= 16'h04DF;
    16'd57668: out <= 16'h0208;    16'd57669: out <= 16'h0211;    16'd57670: out <= 16'h0819;    16'd57671: out <= 16'h01EC;
    16'd57672: out <= 16'h0B0B;    16'd57673: out <= 16'h0624;    16'd57674: out <= 16'h040D;    16'd57675: out <= 16'h0208;
    16'd57676: out <= 16'h043F;    16'd57677: out <= 16'h0462;    16'd57678: out <= 16'h0839;    16'd57679: out <= 16'h06A5;
    16'd57680: out <= 16'h0166;    16'd57681: out <= 16'h056F;    16'd57682: out <= 16'h0301;    16'd57683: out <= 16'h02A4;
    16'd57684: out <= 16'h04BA;    16'd57685: out <= 16'h038C;    16'd57686: out <= 16'h0537;    16'd57687: out <= 16'h0109;
    16'd57688: out <= 16'h0889;    16'd57689: out <= 16'h09FD;    16'd57690: out <= 16'h03CC;    16'd57691: out <= 16'h07B9;
    16'd57692: out <= 16'h0001;    16'd57693: out <= 16'h0236;    16'd57694: out <= 16'h05ED;    16'd57695: out <= 16'h0735;
    16'd57696: out <= 16'h04A0;    16'd57697: out <= 16'h059E;    16'd57698: out <= 16'h0551;    16'd57699: out <= 16'hFF53;
    16'd57700: out <= 16'h0705;    16'd57701: out <= 16'h0933;    16'd57702: out <= 16'h04E3;    16'd57703: out <= 16'h03D7;
    16'd57704: out <= 16'h0128;    16'd57705: out <= 16'hFDA9;    16'd57706: out <= 16'h017F;    16'd57707: out <= 16'h09C9;
    16'd57708: out <= 16'h0478;    16'd57709: out <= 16'h011F;    16'd57710: out <= 16'h00AB;    16'd57711: out <= 16'h04F2;
    16'd57712: out <= 16'h0773;    16'd57713: out <= 16'h06BF;    16'd57714: out <= 16'h075A;    16'd57715: out <= 16'h0659;
    16'd57716: out <= 16'h02C6;    16'd57717: out <= 16'h055D;    16'd57718: out <= 16'h0428;    16'd57719: out <= 16'h0746;
    16'd57720: out <= 16'hFEBA;    16'd57721: out <= 16'h032F;    16'd57722: out <= 16'h0656;    16'd57723: out <= 16'h032F;
    16'd57724: out <= 16'h0373;    16'd57725: out <= 16'h00F1;    16'd57726: out <= 16'h0061;    16'd57727: out <= 16'hFEFC;
    16'd57728: out <= 16'h065F;    16'd57729: out <= 16'h040F;    16'd57730: out <= 16'h0325;    16'd57731: out <= 16'h029B;
    16'd57732: out <= 16'h086A;    16'd57733: out <= 16'hFF73;    16'd57734: out <= 16'hFE21;    16'd57735: out <= 16'hFFCE;
    16'd57736: out <= 16'h03F5;    16'd57737: out <= 16'h06D5;    16'd57738: out <= 16'h0440;    16'd57739: out <= 16'h051C;
    16'd57740: out <= 16'h0890;    16'd57741: out <= 16'h05A4;    16'd57742: out <= 16'h0309;    16'd57743: out <= 16'hFB07;
    16'd57744: out <= 16'h0830;    16'd57745: out <= 16'h079D;    16'd57746: out <= 16'h0846;    16'd57747: out <= 16'hFC98;
    16'd57748: out <= 16'h00A9;    16'd57749: out <= 16'h0222;    16'd57750: out <= 16'h040E;    16'd57751: out <= 16'h02A4;
    16'd57752: out <= 16'h0399;    16'd57753: out <= 16'h0313;    16'd57754: out <= 16'h0719;    16'd57755: out <= 16'h07A4;
    16'd57756: out <= 16'h0225;    16'd57757: out <= 16'h03DD;    16'd57758: out <= 16'hFE75;    16'd57759: out <= 16'h03A7;
    16'd57760: out <= 16'h048D;    16'd57761: out <= 16'h0517;    16'd57762: out <= 16'h0473;    16'd57763: out <= 16'h0324;
    16'd57764: out <= 16'h092C;    16'd57765: out <= 16'h03C4;    16'd57766: out <= 16'h0342;    16'd57767: out <= 16'h05D5;
    16'd57768: out <= 16'h0B5A;    16'd57769: out <= 16'h0612;    16'd57770: out <= 16'h0692;    16'd57771: out <= 16'h019A;
    16'd57772: out <= 16'h0798;    16'd57773: out <= 16'h0066;    16'd57774: out <= 16'h0096;    16'd57775: out <= 16'h0472;
    16'd57776: out <= 16'hFD31;    16'd57777: out <= 16'h052F;    16'd57778: out <= 16'h03A1;    16'd57779: out <= 16'hFD94;
    16'd57780: out <= 16'h0814;    16'd57781: out <= 16'h02B3;    16'd57782: out <= 16'h03CC;    16'd57783: out <= 16'h053A;
    16'd57784: out <= 16'hFCE0;    16'd57785: out <= 16'h0023;    16'd57786: out <= 16'h04D8;    16'd57787: out <= 16'h0B20;
    16'd57788: out <= 16'h0BDB;    16'd57789: out <= 16'h04EF;    16'd57790: out <= 16'h02CB;    16'd57791: out <= 16'h0219;
    16'd57792: out <= 16'h0548;    16'd57793: out <= 16'h01F3;    16'd57794: out <= 16'h0321;    16'd57795: out <= 16'h0279;
    16'd57796: out <= 16'hFB1B;    16'd57797: out <= 16'hFDF8;    16'd57798: out <= 16'h06D0;    16'd57799: out <= 16'h0707;
    16'd57800: out <= 16'h01CE;    16'd57801: out <= 16'h0279;    16'd57802: out <= 16'hFC42;    16'd57803: out <= 16'hFA13;
    16'd57804: out <= 16'hFDBC;    16'd57805: out <= 16'hFEED;    16'd57806: out <= 16'h0058;    16'd57807: out <= 16'h05AF;
    16'd57808: out <= 16'hFE17;    16'd57809: out <= 16'h007E;    16'd57810: out <= 16'h00C6;    16'd57811: out <= 16'hFF61;
    16'd57812: out <= 16'h024C;    16'd57813: out <= 16'h0638;    16'd57814: out <= 16'h007E;    16'd57815: out <= 16'hFACB;
    16'd57816: out <= 16'h02C9;    16'd57817: out <= 16'h01AF;    16'd57818: out <= 16'hFF2C;    16'd57819: out <= 16'h0237;
    16'd57820: out <= 16'hFDD0;    16'd57821: out <= 16'h0179;    16'd57822: out <= 16'hFCE7;    16'd57823: out <= 16'h0193;
    16'd57824: out <= 16'h0135;    16'd57825: out <= 16'hFE3F;    16'd57826: out <= 16'h000A;    16'd57827: out <= 16'h0062;
    16'd57828: out <= 16'hFCD5;    16'd57829: out <= 16'h01B6;    16'd57830: out <= 16'hFBB2;    16'd57831: out <= 16'h0004;
    16'd57832: out <= 16'h027D;    16'd57833: out <= 16'hFE56;    16'd57834: out <= 16'h027E;    16'd57835: out <= 16'hFE23;
    16'd57836: out <= 16'hF847;    16'd57837: out <= 16'hFB33;    16'd57838: out <= 16'hFCBC;    16'd57839: out <= 16'h05EC;
    16'd57840: out <= 16'hF5DE;    16'd57841: out <= 16'hFAAE;    16'd57842: out <= 16'hFC7C;    16'd57843: out <= 16'hFFA2;
    16'd57844: out <= 16'h02BA;    16'd57845: out <= 16'hFBCE;    16'd57846: out <= 16'h0271;    16'd57847: out <= 16'h02A3;
    16'd57848: out <= 16'h02C8;    16'd57849: out <= 16'h045D;    16'd57850: out <= 16'h015D;    16'd57851: out <= 16'hFF2F;
    16'd57852: out <= 16'hFEAF;    16'd57853: out <= 16'h0177;    16'd57854: out <= 16'hFB59;    16'd57855: out <= 16'hFFD3;
    16'd57856: out <= 16'hFCBC;    16'd57857: out <= 16'h02AA;    16'd57858: out <= 16'h01DD;    16'd57859: out <= 16'h0032;
    16'd57860: out <= 16'hFFF3;    16'd57861: out <= 16'hFA01;    16'd57862: out <= 16'h009D;    16'd57863: out <= 16'h0461;
    16'd57864: out <= 16'hFEC2;    16'd57865: out <= 16'h05C6;    16'd57866: out <= 16'h00BC;    16'd57867: out <= 16'h014D;
    16'd57868: out <= 16'hFF67;    16'd57869: out <= 16'h0388;    16'd57870: out <= 16'h05BA;    16'd57871: out <= 16'hFECE;
    16'd57872: out <= 16'hFB3F;    16'd57873: out <= 16'hFBD7;    16'd57874: out <= 16'h01A6;    16'd57875: out <= 16'hFF69;
    16'd57876: out <= 16'h007B;    16'd57877: out <= 16'hFADF;    16'd57878: out <= 16'h008C;    16'd57879: out <= 16'hF9A3;
    16'd57880: out <= 16'h017B;    16'd57881: out <= 16'h03B2;    16'd57882: out <= 16'hFD29;    16'd57883: out <= 16'hFE99;
    16'd57884: out <= 16'hFDFB;    16'd57885: out <= 16'hF7F5;    16'd57886: out <= 16'h04FE;    16'd57887: out <= 16'hFC85;
    16'd57888: out <= 16'hFE20;    16'd57889: out <= 16'hFEC6;    16'd57890: out <= 16'hFFF4;    16'd57891: out <= 16'hF9BE;
    16'd57892: out <= 16'h0721;    16'd57893: out <= 16'hFFCF;    16'd57894: out <= 16'hFFEF;    16'd57895: out <= 16'h037A;
    16'd57896: out <= 16'hFFAD;    16'd57897: out <= 16'h03AD;    16'd57898: out <= 16'hFD7B;    16'd57899: out <= 16'h0538;
    16'd57900: out <= 16'h007F;    16'd57901: out <= 16'hFDE0;    16'd57902: out <= 16'hF832;    16'd57903: out <= 16'hFFD8;
    16'd57904: out <= 16'h0543;    16'd57905: out <= 16'h03CB;    16'd57906: out <= 16'h0560;    16'd57907: out <= 16'h01CC;
    16'd57908: out <= 16'h07FF;    16'd57909: out <= 16'h05F6;    16'd57910: out <= 16'h048B;    16'd57911: out <= 16'h03CC;
    16'd57912: out <= 16'hFE9D;    16'd57913: out <= 16'h00C8;    16'd57914: out <= 16'hFAAD;    16'd57915: out <= 16'h03D3;
    16'd57916: out <= 16'h019B;    16'd57917: out <= 16'h03BB;    16'd57918: out <= 16'h07CD;    16'd57919: out <= 16'h0714;
    16'd57920: out <= 16'h02BD;    16'd57921: out <= 16'h047A;    16'd57922: out <= 16'h05F5;    16'd57923: out <= 16'h0476;
    16'd57924: out <= 16'h0051;    16'd57925: out <= 16'h001E;    16'd57926: out <= 16'h02AC;    16'd57927: out <= 16'h05CF;
    16'd57928: out <= 16'h034A;    16'd57929: out <= 16'h02AB;    16'd57930: out <= 16'h061E;    16'd57931: out <= 16'h0036;
    16'd57932: out <= 16'hFA47;    16'd57933: out <= 16'h054B;    16'd57934: out <= 16'h058B;    16'd57935: out <= 16'hFD32;
    16'd57936: out <= 16'h0288;    16'd57937: out <= 16'h0309;    16'd57938: out <= 16'h05DE;    16'd57939: out <= 16'h0672;
    16'd57940: out <= 16'h055D;    16'd57941: out <= 16'hFEE3;    16'd57942: out <= 16'h06BD;    16'd57943: out <= 16'h0390;
    16'd57944: out <= 16'h028F;    16'd57945: out <= 16'h0923;    16'd57946: out <= 16'h0752;    16'd57947: out <= 16'h084D;
    16'd57948: out <= 16'h081C;    16'd57949: out <= 16'h07AF;    16'd57950: out <= 16'h016A;    16'd57951: out <= 16'h0989;
    16'd57952: out <= 16'h0082;    16'd57953: out <= 16'h0357;    16'd57954: out <= 16'h0018;    16'd57955: out <= 16'h029F;
    16'd57956: out <= 16'h01CB;    16'd57957: out <= 16'h04D0;    16'd57958: out <= 16'h0580;    16'd57959: out <= 16'hFF7F;
    16'd57960: out <= 16'h04D8;    16'd57961: out <= 16'h0770;    16'd57962: out <= 16'h0849;    16'd57963: out <= 16'h00C6;
    16'd57964: out <= 16'h0099;    16'd57965: out <= 16'h0131;    16'd57966: out <= 16'h06A6;    16'd57967: out <= 16'h0873;
    16'd57968: out <= 16'hFEEC;    16'd57969: out <= 16'hFF0B;    16'd57970: out <= 16'h0B3B;    16'd57971: out <= 16'h06D1;
    16'd57972: out <= 16'h02BB;    16'd57973: out <= 16'h0292;    16'd57974: out <= 16'h09FE;    16'd57975: out <= 16'h051D;
    16'd57976: out <= 16'h04E5;    16'd57977: out <= 16'h0202;    16'd57978: out <= 16'h0AAB;    16'd57979: out <= 16'h0302;
    16'd57980: out <= 16'hFF4B;    16'd57981: out <= 16'h0468;    16'd57982: out <= 16'h0066;    16'd57983: out <= 16'hFFF7;
    16'd57984: out <= 16'h092A;    16'd57985: out <= 16'h048E;    16'd57986: out <= 16'h005F;    16'd57987: out <= 16'h0060;
    16'd57988: out <= 16'hF8CA;    16'd57989: out <= 16'h0792;    16'd57990: out <= 16'h0453;    16'd57991: out <= 16'h030D;
    16'd57992: out <= 16'h054E;    16'd57993: out <= 16'h015F;    16'd57994: out <= 16'h0330;    16'd57995: out <= 16'h0835;
    16'd57996: out <= 16'h0297;    16'd57997: out <= 16'h011F;    16'd57998: out <= 16'h00D8;    16'd57999: out <= 16'hFDA6;
    16'd58000: out <= 16'h0901;    16'd58001: out <= 16'hFC6A;    16'd58002: out <= 16'h0796;    16'd58003: out <= 16'hFF6C;
    16'd58004: out <= 16'h06D4;    16'd58005: out <= 16'h04EB;    16'd58006: out <= 16'h0CD7;    16'd58007: out <= 16'h03C5;
    16'd58008: out <= 16'h0234;    16'd58009: out <= 16'h01CA;    16'd58010: out <= 16'h0673;    16'd58011: out <= 16'h0477;
    16'd58012: out <= 16'hFF8A;    16'd58013: out <= 16'h01C6;    16'd58014: out <= 16'h02BA;    16'd58015: out <= 16'h02F4;
    16'd58016: out <= 16'h0335;    16'd58017: out <= 16'hFBEB;    16'd58018: out <= 16'h09A8;    16'd58019: out <= 16'h022E;
    16'd58020: out <= 16'h0385;    16'd58021: out <= 16'h0145;    16'd58022: out <= 16'h003B;    16'd58023: out <= 16'h006E;
    16'd58024: out <= 16'hFEBA;    16'd58025: out <= 16'h0638;    16'd58026: out <= 16'h057E;    16'd58027: out <= 16'h0015;
    16'd58028: out <= 16'hFCD6;    16'd58029: out <= 16'h075A;    16'd58030: out <= 16'h05B3;    16'd58031: out <= 16'hFD15;
    16'd58032: out <= 16'h07C5;    16'd58033: out <= 16'h07F8;    16'd58034: out <= 16'hFE38;    16'd58035: out <= 16'h018B;
    16'd58036: out <= 16'h05E4;    16'd58037: out <= 16'hFE54;    16'd58038: out <= 16'h092F;    16'd58039: out <= 16'h007E;
    16'd58040: out <= 16'h08A0;    16'd58041: out <= 16'h0199;    16'd58042: out <= 16'h01ED;    16'd58043: out <= 16'h034E;
    16'd58044: out <= 16'h03FF;    16'd58045: out <= 16'h0378;    16'd58046: out <= 16'h0C29;    16'd58047: out <= 16'h0230;
    16'd58048: out <= 16'h028B;    16'd58049: out <= 16'hFFC2;    16'd58050: out <= 16'hFBF1;    16'd58051: out <= 16'hFDB4;
    16'd58052: out <= 16'hFF91;    16'd58053: out <= 16'h06A1;    16'd58054: out <= 16'h054F;    16'd58055: out <= 16'h0187;
    16'd58056: out <= 16'hFD05;    16'd58057: out <= 16'h0514;    16'd58058: out <= 16'h06F5;    16'd58059: out <= 16'hF895;
    16'd58060: out <= 16'h018E;    16'd58061: out <= 16'hF869;    16'd58062: out <= 16'h0000;    16'd58063: out <= 16'hF9F6;
    16'd58064: out <= 16'hFBC1;    16'd58065: out <= 16'h02E2;    16'd58066: out <= 16'hFAEF;    16'd58067: out <= 16'h014B;
    16'd58068: out <= 16'h00CD;    16'd58069: out <= 16'h0462;    16'd58070: out <= 16'hFE7D;    16'd58071: out <= 16'hFCC6;
    16'd58072: out <= 16'h08D6;    16'd58073: out <= 16'h0413;    16'd58074: out <= 16'h0500;    16'd58075: out <= 16'h048D;
    16'd58076: out <= 16'hFC03;    16'd58077: out <= 16'hFD60;    16'd58078: out <= 16'hFD44;    16'd58079: out <= 16'hFC4C;
    16'd58080: out <= 16'hF6B1;    16'd58081: out <= 16'hFDFE;    16'd58082: out <= 16'h04D2;    16'd58083: out <= 16'h0020;
    16'd58084: out <= 16'h011C;    16'd58085: out <= 16'h001B;    16'd58086: out <= 16'h0280;    16'd58087: out <= 16'hFABB;
    16'd58088: out <= 16'h0287;    16'd58089: out <= 16'hFC3B;    16'd58090: out <= 16'hF867;    16'd58091: out <= 16'h02FD;
    16'd58092: out <= 16'hFF4D;    16'd58093: out <= 16'h02B4;    16'd58094: out <= 16'hFF4A;    16'd58095: out <= 16'hFFDF;
    16'd58096: out <= 16'h0235;    16'd58097: out <= 16'hFF1D;    16'd58098: out <= 16'hFDC3;    16'd58099: out <= 16'hFC0F;
    16'd58100: out <= 16'h03B8;    16'd58101: out <= 16'h03D0;    16'd58102: out <= 16'h01DF;    16'd58103: out <= 16'h05A6;
    16'd58104: out <= 16'h01E9;    16'd58105: out <= 16'hFAF4;    16'd58106: out <= 16'h0098;    16'd58107: out <= 16'hFF0A;
    16'd58108: out <= 16'h0611;    16'd58109: out <= 16'h00F1;    16'd58110: out <= 16'h0442;    16'd58111: out <= 16'h02E0;
    16'd58112: out <= 16'h00C9;    16'd58113: out <= 16'hFD94;    16'd58114: out <= 16'hF887;    16'd58115: out <= 16'h03DB;
    16'd58116: out <= 16'h0076;    16'd58117: out <= 16'hFF5E;    16'd58118: out <= 16'hFC84;    16'd58119: out <= 16'hF975;
    16'd58120: out <= 16'hF92E;    16'd58121: out <= 16'h00EC;    16'd58122: out <= 16'h0054;    16'd58123: out <= 16'hF88D;
    16'd58124: out <= 16'h05BC;    16'd58125: out <= 16'hFA24;    16'd58126: out <= 16'h04B1;    16'd58127: out <= 16'h0284;
    16'd58128: out <= 16'h0133;    16'd58129: out <= 16'hFD10;    16'd58130: out <= 16'hFBA0;    16'd58131: out <= 16'h0752;
    16'd58132: out <= 16'h010F;    16'd58133: out <= 16'h0698;    16'd58134: out <= 16'h02F5;    16'd58135: out <= 16'hFE01;
    16'd58136: out <= 16'hFBE2;    16'd58137: out <= 16'hFDCB;    16'd58138: out <= 16'h008D;    16'd58139: out <= 16'h02FF;
    16'd58140: out <= 16'hFF2A;    16'd58141: out <= 16'hFD06;    16'd58142: out <= 16'hFFCA;    16'd58143: out <= 16'h0576;
    16'd58144: out <= 16'hFB9D;    16'd58145: out <= 16'h059D;    16'd58146: out <= 16'h0357;    16'd58147: out <= 16'h060D;
    16'd58148: out <= 16'hFD81;    16'd58149: out <= 16'hFB9E;    16'd58150: out <= 16'h010E;    16'd58151: out <= 16'hFE61;
    16'd58152: out <= 16'h06E9;    16'd58153: out <= 16'hFD43;    16'd58154: out <= 16'hFA56;    16'd58155: out <= 16'hFB63;
    16'd58156: out <= 16'hFFA5;    16'd58157: out <= 16'hFCDA;    16'd58158: out <= 16'h0037;    16'd58159: out <= 16'h038B;
    16'd58160: out <= 16'hFF0C;    16'd58161: out <= 16'h0917;    16'd58162: out <= 16'h0234;    16'd58163: out <= 16'h0C67;
    16'd58164: out <= 16'h0610;    16'd58165: out <= 16'h037D;    16'd58166: out <= 16'h0BD4;    16'd58167: out <= 16'h01AA;
    16'd58168: out <= 16'h0474;    16'd58169: out <= 16'h028D;    16'd58170: out <= 16'h086C;    16'd58171: out <= 16'h0358;
    16'd58172: out <= 16'h05A9;    16'd58173: out <= 16'hFFF3;    16'd58174: out <= 16'h000E;    16'd58175: out <= 16'h08FE;
    16'd58176: out <= 16'h0208;    16'd58177: out <= 16'h065F;    16'd58178: out <= 16'h0669;    16'd58179: out <= 16'h0D40;
    16'd58180: out <= 16'h00B5;    16'd58181: out <= 16'h037C;    16'd58182: out <= 16'h07E5;    16'd58183: out <= 16'h0317;
    16'd58184: out <= 16'h096E;    16'd58185: out <= 16'h0953;    16'd58186: out <= 16'h0B54;    16'd58187: out <= 16'h04B1;
    16'd58188: out <= 16'h0787;    16'd58189: out <= 16'h03A8;    16'd58190: out <= 16'h06C6;    16'd58191: out <= 16'h07D1;
    16'd58192: out <= 16'h02AF;    16'd58193: out <= 16'h05FC;    16'd58194: out <= 16'h0762;    16'd58195: out <= 16'hFE49;
    16'd58196: out <= 16'h0875;    16'd58197: out <= 16'hFFB0;    16'd58198: out <= 16'hF99B;    16'd58199: out <= 16'h025A;
    16'd58200: out <= 16'h02D8;    16'd58201: out <= 16'h06E8;    16'd58202: out <= 16'hFFCE;    16'd58203: out <= 16'h07BE;
    16'd58204: out <= 16'hFFB5;    16'd58205: out <= 16'hFCF2;    16'd58206: out <= 16'h0452;    16'd58207: out <= 16'h0A15;
    16'd58208: out <= 16'h0356;    16'd58209: out <= 16'h05E9;    16'd58210: out <= 16'hFFC5;    16'd58211: out <= 16'h00A5;
    16'd58212: out <= 16'h03E4;    16'd58213: out <= 16'h0797;    16'd58214: out <= 16'h0400;    16'd58215: out <= 16'h055A;
    16'd58216: out <= 16'hFBDE;    16'd58217: out <= 16'h086D;    16'd58218: out <= 16'hFF42;    16'd58219: out <= 16'hFF22;
    16'd58220: out <= 16'h0220;    16'd58221: out <= 16'hFA95;    16'd58222: out <= 16'h082E;    16'd58223: out <= 16'h05D1;
    16'd58224: out <= 16'h04EE;    16'd58225: out <= 16'h01F2;    16'd58226: out <= 16'hFFDD;    16'd58227: out <= 16'h038C;
    16'd58228: out <= 16'hFFE5;    16'd58229: out <= 16'h0390;    16'd58230: out <= 16'h06D0;    16'd58231: out <= 16'hFFFC;
    16'd58232: out <= 16'h0B81;    16'd58233: out <= 16'hFF82;    16'd58234: out <= 16'h0380;    16'd58235: out <= 16'hFFB0;
    16'd58236: out <= 16'h0883;    16'd58237: out <= 16'h053D;    16'd58238: out <= 16'h0209;    16'd58239: out <= 16'h0447;
    16'd58240: out <= 16'hFFC3;    16'd58241: out <= 16'h020E;    16'd58242: out <= 16'h006E;    16'd58243: out <= 16'h05D9;
    16'd58244: out <= 16'hFDBA;    16'd58245: out <= 16'h0918;    16'd58246: out <= 16'h0682;    16'd58247: out <= 16'h02F1;
    16'd58248: out <= 16'hFC73;    16'd58249: out <= 16'h05BB;    16'd58250: out <= 16'hFE13;    16'd58251: out <= 16'h00A9;
    16'd58252: out <= 16'hFD77;    16'd58253: out <= 16'h0C48;    16'd58254: out <= 16'h0511;    16'd58255: out <= 16'h028D;
    16'd58256: out <= 16'h067D;    16'd58257: out <= 16'hFE0F;    16'd58258: out <= 16'h05CE;    16'd58259: out <= 16'hFF5B;
    16'd58260: out <= 16'h05A0;    16'd58261: out <= 16'hFF55;    16'd58262: out <= 16'hFCE0;    16'd58263: out <= 16'h0667;
    16'd58264: out <= 16'h06CE;    16'd58265: out <= 16'h010F;    16'd58266: out <= 16'h024F;    16'd58267: out <= 16'hFDB6;
    16'd58268: out <= 16'h0547;    16'd58269: out <= 16'h01AB;    16'd58270: out <= 16'h0B4F;    16'd58271: out <= 16'hFA83;
    16'd58272: out <= 16'h05F1;    16'd58273: out <= 16'h0455;    16'd58274: out <= 16'hFD3F;    16'd58275: out <= 16'h030E;
    16'd58276: out <= 16'hFE6F;    16'd58277: out <= 16'h01C8;    16'd58278: out <= 16'h09AE;    16'd58279: out <= 16'h0A3E;
    16'd58280: out <= 16'h02AA;    16'd58281: out <= 16'h0174;    16'd58282: out <= 16'h0397;    16'd58283: out <= 16'h02FB;
    16'd58284: out <= 16'h017A;    16'd58285: out <= 16'h0122;    16'd58286: out <= 16'hFCBF;    16'd58287: out <= 16'h0015;
    16'd58288: out <= 16'h0531;    16'd58289: out <= 16'h032D;    16'd58290: out <= 16'h0746;    16'd58291: out <= 16'h06D4;
    16'd58292: out <= 16'h0524;    16'd58293: out <= 16'h00BA;    16'd58294: out <= 16'hFCF4;    16'd58295: out <= 16'h0B03;
    16'd58296: out <= 16'h0272;    16'd58297: out <= 16'hFE9F;    16'd58298: out <= 16'h0275;    16'd58299: out <= 16'h01A3;
    16'd58300: out <= 16'hFE6F;    16'd58301: out <= 16'h0248;    16'd58302: out <= 16'h06AE;    16'd58303: out <= 16'h04A8;
    16'd58304: out <= 16'h08A5;    16'd58305: out <= 16'h0151;    16'd58306: out <= 16'h08A1;    16'd58307: out <= 16'h01CB;
    16'd58308: out <= 16'hFE66;    16'd58309: out <= 16'hFE27;    16'd58310: out <= 16'hFE36;    16'd58311: out <= 16'hFBC9;
    16'd58312: out <= 16'h02C3;    16'd58313: out <= 16'hFE12;    16'd58314: out <= 16'hFB59;    16'd58315: out <= 16'hF714;
    16'd58316: out <= 16'h0373;    16'd58317: out <= 16'hFE57;    16'd58318: out <= 16'hFF94;    16'd58319: out <= 16'h0A51;
    16'd58320: out <= 16'h00CE;    16'd58321: out <= 16'h0000;    16'd58322: out <= 16'h02DE;    16'd58323: out <= 16'h04AD;
    16'd58324: out <= 16'h0171;    16'd58325: out <= 16'hFE41;    16'd58326: out <= 16'hFD6A;    16'd58327: out <= 16'h01F9;
    16'd58328: out <= 16'h02F9;    16'd58329: out <= 16'hFD13;    16'd58330: out <= 16'hF981;    16'd58331: out <= 16'hFF20;
    16'd58332: out <= 16'h008B;    16'd58333: out <= 16'h0464;    16'd58334: out <= 16'h0B79;    16'd58335: out <= 16'h01AB;
    16'd58336: out <= 16'hFCEE;    16'd58337: out <= 16'h037F;    16'd58338: out <= 16'hFCD7;    16'd58339: out <= 16'hFBB7;
    16'd58340: out <= 16'h03CD;    16'd58341: out <= 16'h0148;    16'd58342: out <= 16'h00AA;    16'd58343: out <= 16'hF9F0;
    16'd58344: out <= 16'h0045;    16'd58345: out <= 16'hFEB6;    16'd58346: out <= 16'h025B;    16'd58347: out <= 16'hFF86;
    16'd58348: out <= 16'hFEFE;    16'd58349: out <= 16'h01CA;    16'd58350: out <= 16'h032A;    16'd58351: out <= 16'h0049;
    16'd58352: out <= 16'hFEE6;    16'd58353: out <= 16'h04DA;    16'd58354: out <= 16'hFB3B;    16'd58355: out <= 16'h0285;
    16'd58356: out <= 16'h065E;    16'd58357: out <= 16'hFEAD;    16'd58358: out <= 16'h03E6;    16'd58359: out <= 16'h024A;
    16'd58360: out <= 16'hFDED;    16'd58361: out <= 16'h0188;    16'd58362: out <= 16'hFDE1;    16'd58363: out <= 16'hFB2C;
    16'd58364: out <= 16'h04CC;    16'd58365: out <= 16'hFFE6;    16'd58366: out <= 16'h03B9;    16'd58367: out <= 16'h00E0;
    16'd58368: out <= 16'hFF4B;    16'd58369: out <= 16'hFC7D;    16'd58370: out <= 16'h00EC;    16'd58371: out <= 16'h022C;
    16'd58372: out <= 16'hF5EB;    16'd58373: out <= 16'hFE4F;    16'd58374: out <= 16'h0551;    16'd58375: out <= 16'hFC12;
    16'd58376: out <= 16'hFE84;    16'd58377: out <= 16'h004D;    16'd58378: out <= 16'hFA44;    16'd58379: out <= 16'h032C;
    16'd58380: out <= 16'hF83D;    16'd58381: out <= 16'hFB75;    16'd58382: out <= 16'hFE8D;    16'd58383: out <= 16'hF90C;
    16'd58384: out <= 16'hFBAD;    16'd58385: out <= 16'hFFAC;    16'd58386: out <= 16'h035A;    16'd58387: out <= 16'h0248;
    16'd58388: out <= 16'h02AB;    16'd58389: out <= 16'h0848;    16'd58390: out <= 16'hFB3A;    16'd58391: out <= 16'hFD08;
    16'd58392: out <= 16'hFC7A;    16'd58393: out <= 16'hFFEF;    16'd58394: out <= 16'h00E4;    16'd58395: out <= 16'hFF9E;
    16'd58396: out <= 16'h02C4;    16'd58397: out <= 16'hFE56;    16'd58398: out <= 16'h0860;    16'd58399: out <= 16'hFDBF;
    16'd58400: out <= 16'hFD1E;    16'd58401: out <= 16'h0095;    16'd58402: out <= 16'hFE24;    16'd58403: out <= 16'h0469;
    16'd58404: out <= 16'hFD1A;    16'd58405: out <= 16'h002B;    16'd58406: out <= 16'hFEA8;    16'd58407: out <= 16'hFFDD;
    16'd58408: out <= 16'h0368;    16'd58409: out <= 16'hFFCD;    16'd58410: out <= 16'hFB23;    16'd58411: out <= 16'hFD9C;
    16'd58412: out <= 16'h08B3;    16'd58413: out <= 16'h040D;    16'd58414: out <= 16'hFBFC;    16'd58415: out <= 16'h0091;
    16'd58416: out <= 16'h0739;    16'd58417: out <= 16'h0826;    16'd58418: out <= 16'h0112;    16'd58419: out <= 16'h0532;
    16'd58420: out <= 16'h00AA;    16'd58421: out <= 16'h0537;    16'd58422: out <= 16'h0360;    16'd58423: out <= 16'h00FC;
    16'd58424: out <= 16'h0631;    16'd58425: out <= 16'hFD9D;    16'd58426: out <= 16'hFE57;    16'd58427: out <= 16'h022F;
    16'd58428: out <= 16'h02ED;    16'd58429: out <= 16'h05CF;    16'd58430: out <= 16'h06F3;    16'd58431: out <= 16'h01A9;
    16'd58432: out <= 16'h0808;    16'd58433: out <= 16'h06CB;    16'd58434: out <= 16'hFF5C;    16'd58435: out <= 16'h098C;
    16'd58436: out <= 16'h05C1;    16'd58437: out <= 16'hFF98;    16'd58438: out <= 16'h0166;    16'd58439: out <= 16'h0675;
    16'd58440: out <= 16'h01C5;    16'd58441: out <= 16'h0425;    16'd58442: out <= 16'h012B;    16'd58443: out <= 16'h062B;
    16'd58444: out <= 16'h0634;    16'd58445: out <= 16'h00B6;    16'd58446: out <= 16'h09AA;    16'd58447: out <= 16'h081B;
    16'd58448: out <= 16'h0302;    16'd58449: out <= 16'h059E;    16'd58450: out <= 16'h05A3;    16'd58451: out <= 16'h074E;
    16'd58452: out <= 16'h0495;    16'd58453: out <= 16'hFF4E;    16'd58454: out <= 16'h07D2;    16'd58455: out <= 16'h0417;
    16'd58456: out <= 16'h008B;    16'd58457: out <= 16'h0674;    16'd58458: out <= 16'hFD45;    16'd58459: out <= 16'h06BE;
    16'd58460: out <= 16'h06F0;    16'd58461: out <= 16'h00BC;    16'd58462: out <= 16'h03D8;    16'd58463: out <= 16'h0550;
    16'd58464: out <= 16'h07D4;    16'd58465: out <= 16'h0633;    16'd58466: out <= 16'h05A1;    16'd58467: out <= 16'h0246;
    16'd58468: out <= 16'h022E;    16'd58469: out <= 16'h03DE;    16'd58470: out <= 16'h0121;    16'd58471: out <= 16'h04AF;
    16'd58472: out <= 16'h0156;    16'd58473: out <= 16'hFE5C;    16'd58474: out <= 16'h0210;    16'd58475: out <= 16'h00DC;
    16'd58476: out <= 16'h016F;    16'd58477: out <= 16'h08CD;    16'd58478: out <= 16'h0351;    16'd58479: out <= 16'h0C17;
    16'd58480: out <= 16'h0624;    16'd58481: out <= 16'h0094;    16'd58482: out <= 16'h0560;    16'd58483: out <= 16'h04E1;
    16'd58484: out <= 16'h049D;    16'd58485: out <= 16'h04D4;    16'd58486: out <= 16'h0815;    16'd58487: out <= 16'h00A1;
    16'd58488: out <= 16'h0755;    16'd58489: out <= 16'hFD5E;    16'd58490: out <= 16'h072B;    16'd58491: out <= 16'h05DA;
    16'd58492: out <= 16'h051B;    16'd58493: out <= 16'hFEE8;    16'd58494: out <= 16'h080C;    16'd58495: out <= 16'h02B6;
    16'd58496: out <= 16'hFE73;    16'd58497: out <= 16'h08E5;    16'd58498: out <= 16'h041F;    16'd58499: out <= 16'h0415;
    16'd58500: out <= 16'h052F;    16'd58501: out <= 16'h016D;    16'd58502: out <= 16'h0857;    16'd58503: out <= 16'hFCE5;
    16'd58504: out <= 16'h03EA;    16'd58505: out <= 16'hFECE;    16'd58506: out <= 16'h0515;    16'd58507: out <= 16'h023B;
    16'd58508: out <= 16'h05E8;    16'd58509: out <= 16'h00DA;    16'd58510: out <= 16'h0248;    16'd58511: out <= 16'h0367;
    16'd58512: out <= 16'hFDCF;    16'd58513: out <= 16'h0560;    16'd58514: out <= 16'h0328;    16'd58515: out <= 16'h030D;
    16'd58516: out <= 16'hFA7D;    16'd58517: out <= 16'h004F;    16'd58518: out <= 16'hFCD0;    16'd58519: out <= 16'h098A;
    16'd58520: out <= 16'hFF5D;    16'd58521: out <= 16'h0593;    16'd58522: out <= 16'h08C0;    16'd58523: out <= 16'hFEB9;
    16'd58524: out <= 16'h01CE;    16'd58525: out <= 16'h049E;    16'd58526: out <= 16'h0A30;    16'd58527: out <= 16'h04F6;
    16'd58528: out <= 16'h0305;    16'd58529: out <= 16'h0528;    16'd58530: out <= 16'h06D5;    16'd58531: out <= 16'h048C;
    16'd58532: out <= 16'hFEB8;    16'd58533: out <= 16'h0448;    16'd58534: out <= 16'h0AD0;    16'd58535: out <= 16'h07EE;
    16'd58536: out <= 16'h00EA;    16'd58537: out <= 16'h0264;    16'd58538: out <= 16'h0625;    16'd58539: out <= 16'h0945;
    16'd58540: out <= 16'hFC19;    16'd58541: out <= 16'h04F0;    16'd58542: out <= 16'hFCB4;    16'd58543: out <= 16'h036C;
    16'd58544: out <= 16'h08E8;    16'd58545: out <= 16'hFD8D;    16'd58546: out <= 16'hFCCE;    16'd58547: out <= 16'h0272;
    16'd58548: out <= 16'h085B;    16'd58549: out <= 16'h0784;    16'd58550: out <= 16'h0B04;    16'd58551: out <= 16'hFDDE;
    16'd58552: out <= 16'h03DE;    16'd58553: out <= 16'h061B;    16'd58554: out <= 16'hFEA7;    16'd58555: out <= 16'h044D;
    16'd58556: out <= 16'hFF1B;    16'd58557: out <= 16'h00F0;    16'd58558: out <= 16'h05EB;    16'd58559: out <= 16'h00FF;
    16'd58560: out <= 16'h047B;    16'd58561: out <= 16'h0772;    16'd58562: out <= 16'h08AA;    16'd58563: out <= 16'h01BA;
    16'd58564: out <= 16'h0037;    16'd58565: out <= 16'hFD0D;    16'd58566: out <= 16'h01A6;    16'd58567: out <= 16'hFD5A;
    16'd58568: out <= 16'hFCA0;    16'd58569: out <= 16'hFB5F;    16'd58570: out <= 16'hFF97;    16'd58571: out <= 16'h021E;
    16'd58572: out <= 16'hFFB1;    16'd58573: out <= 16'hFAB4;    16'd58574: out <= 16'h01FA;    16'd58575: out <= 16'h06B4;
    16'd58576: out <= 16'hF8AA;    16'd58577: out <= 16'h0009;    16'd58578: out <= 16'h009C;    16'd58579: out <= 16'h0727;
    16'd58580: out <= 16'hFD35;    16'd58581: out <= 16'hFDC6;    16'd58582: out <= 16'hF894;    16'd58583: out <= 16'hFEF7;
    16'd58584: out <= 16'h03A5;    16'd58585: out <= 16'hFF74;    16'd58586: out <= 16'hFD4C;    16'd58587: out <= 16'hFED0;
    16'd58588: out <= 16'hFEBB;    16'd58589: out <= 16'hFD01;    16'd58590: out <= 16'hF9E7;    16'd58591: out <= 16'hFFE7;
    16'd58592: out <= 16'h03C3;    16'd58593: out <= 16'h01B1;    16'd58594: out <= 16'h02DF;    16'd58595: out <= 16'hFE45;
    16'd58596: out <= 16'hFE29;    16'd58597: out <= 16'h0739;    16'd58598: out <= 16'h0831;    16'd58599: out <= 16'hFFDD;
    16'd58600: out <= 16'hFE15;    16'd58601: out <= 16'h0165;    16'd58602: out <= 16'hF956;    16'd58603: out <= 16'hFC1F;
    16'd58604: out <= 16'h0480;    16'd58605: out <= 16'h072E;    16'd58606: out <= 16'h02C7;    16'd58607: out <= 16'h06D5;
    16'd58608: out <= 16'h022F;    16'd58609: out <= 16'h0B2F;    16'd58610: out <= 16'hFCA7;    16'd58611: out <= 16'hFD83;
    16'd58612: out <= 16'hFDA2;    16'd58613: out <= 16'hFC1F;    16'd58614: out <= 16'hF883;    16'd58615: out <= 16'h054D;
    16'd58616: out <= 16'hFED1;    16'd58617: out <= 16'h0583;    16'd58618: out <= 16'hFEFB;    16'd58619: out <= 16'h0166;
    16'd58620: out <= 16'hFDA2;    16'd58621: out <= 16'h0520;    16'd58622: out <= 16'hFD8F;    16'd58623: out <= 16'hFBDC;
    16'd58624: out <= 16'hFDBF;    16'd58625: out <= 16'h00CC;    16'd58626: out <= 16'hFB65;    16'd58627: out <= 16'h0290;
    16'd58628: out <= 16'hFF33;    16'd58629: out <= 16'hF838;    16'd58630: out <= 16'hFB4F;    16'd58631: out <= 16'h056E;
    16'd58632: out <= 16'h00B7;    16'd58633: out <= 16'hFF5E;    16'd58634: out <= 16'hFE5E;    16'd58635: out <= 16'h068D;
    16'd58636: out <= 16'h01A0;    16'd58637: out <= 16'hFDAA;    16'd58638: out <= 16'h0656;    16'd58639: out <= 16'h00F2;
    16'd58640: out <= 16'h00CA;    16'd58641: out <= 16'h028B;    16'd58642: out <= 16'h05A4;    16'd58643: out <= 16'h01D3;
    16'd58644: out <= 16'h01ED;    16'd58645: out <= 16'hFDD6;    16'd58646: out <= 16'h0293;    16'd58647: out <= 16'h0027;
    16'd58648: out <= 16'hFFAE;    16'd58649: out <= 16'hFA11;    16'd58650: out <= 16'h00DA;    16'd58651: out <= 16'hFED6;
    16'd58652: out <= 16'h0665;    16'd58653: out <= 16'hF82D;    16'd58654: out <= 16'h01EC;    16'd58655: out <= 16'h06B0;
    16'd58656: out <= 16'h01BB;    16'd58657: out <= 16'hFE41;    16'd58658: out <= 16'hFEB1;    16'd58659: out <= 16'hFD30;
    16'd58660: out <= 16'h0392;    16'd58661: out <= 16'hFFA9;    16'd58662: out <= 16'hFF5F;    16'd58663: out <= 16'h01E7;
    16'd58664: out <= 16'hFEF7;    16'd58665: out <= 16'h0399;    16'd58666: out <= 16'hFF4C;    16'd58667: out <= 16'hFB20;
    16'd58668: out <= 16'h00F7;    16'd58669: out <= 16'h046D;    16'd58670: out <= 16'hFCFA;    16'd58671: out <= 16'h0753;
    16'd58672: out <= 16'h054A;    16'd58673: out <= 16'h062A;    16'd58674: out <= 16'h06E7;    16'd58675: out <= 16'h0735;
    16'd58676: out <= 16'h0631;    16'd58677: out <= 16'h0150;    16'd58678: out <= 16'h03AA;    16'd58679: out <= 16'h0987;
    16'd58680: out <= 16'h0425;    16'd58681: out <= 16'h077B;    16'd58682: out <= 16'h00F9;    16'd58683: out <= 16'h04C2;
    16'd58684: out <= 16'h0880;    16'd58685: out <= 16'h016E;    16'd58686: out <= 16'h0077;    16'd58687: out <= 16'h0126;
    16'd58688: out <= 16'h0769;    16'd58689: out <= 16'h0A76;    16'd58690: out <= 16'h0946;    16'd58691: out <= 16'h0165;
    16'd58692: out <= 16'hFCE9;    16'd58693: out <= 16'h093B;    16'd58694: out <= 16'hFD11;    16'd58695: out <= 16'h05C5;
    16'd58696: out <= 16'h05FD;    16'd58697: out <= 16'h012F;    16'd58698: out <= 16'h0969;    16'd58699: out <= 16'h05C7;
    16'd58700: out <= 16'h0364;    16'd58701: out <= 16'h023D;    16'd58702: out <= 16'h024E;    16'd58703: out <= 16'h047C;
    16'd58704: out <= 16'h0492;    16'd58705: out <= 16'h0831;    16'd58706: out <= 16'h0794;    16'd58707: out <= 16'h077F;
    16'd58708: out <= 16'h0669;    16'd58709: out <= 16'h029D;    16'd58710: out <= 16'h0582;    16'd58711: out <= 16'h0661;
    16'd58712: out <= 16'h097C;    16'd58713: out <= 16'hFDB3;    16'd58714: out <= 16'h01F2;    16'd58715: out <= 16'h052D;
    16'd58716: out <= 16'h03C9;    16'd58717: out <= 16'h067A;    16'd58718: out <= 16'h0444;    16'd58719: out <= 16'h0199;
    16'd58720: out <= 16'h000E;    16'd58721: out <= 16'hFE19;    16'd58722: out <= 16'h0220;    16'd58723: out <= 16'h05C2;
    16'd58724: out <= 16'h0200;    16'd58725: out <= 16'h001A;    16'd58726: out <= 16'h0966;    16'd58727: out <= 16'h036F;
    16'd58728: out <= 16'h0351;    16'd58729: out <= 16'h04EE;    16'd58730: out <= 16'hFEF1;    16'd58731: out <= 16'hFE4F;
    16'd58732: out <= 16'h0276;    16'd58733: out <= 16'h01CA;    16'd58734: out <= 16'h06A3;    16'd58735: out <= 16'hFD24;
    16'd58736: out <= 16'h0320;    16'd58737: out <= 16'h03F7;    16'd58738: out <= 16'h0526;    16'd58739: out <= 16'h070D;
    16'd58740: out <= 16'h040B;    16'd58741: out <= 16'h09AB;    16'd58742: out <= 16'h0CED;    16'd58743: out <= 16'hFD33;
    16'd58744: out <= 16'h01EB;    16'd58745: out <= 16'h0225;    16'd58746: out <= 16'h02CF;    16'd58747: out <= 16'h0372;
    16'd58748: out <= 16'hFE0A;    16'd58749: out <= 16'h03B2;    16'd58750: out <= 16'h06A6;    16'd58751: out <= 16'h0AD8;
    16'd58752: out <= 16'hFED7;    16'd58753: out <= 16'hFDDA;    16'd58754: out <= 16'h04DE;    16'd58755: out <= 16'h05F5;
    16'd58756: out <= 16'hFD4C;    16'd58757: out <= 16'hFEB3;    16'd58758: out <= 16'h0418;    16'd58759: out <= 16'h0289;
    16'd58760: out <= 16'hFA8A;    16'd58761: out <= 16'h0606;    16'd58762: out <= 16'h0673;    16'd58763: out <= 16'h0404;
    16'd58764: out <= 16'h0319;    16'd58765: out <= 16'h07ED;    16'd58766: out <= 16'h060B;    16'd58767: out <= 16'h0685;
    16'd58768: out <= 16'h03D0;    16'd58769: out <= 16'h0871;    16'd58770: out <= 16'h0758;    16'd58771: out <= 16'h043B;
    16'd58772: out <= 16'h0AA1;    16'd58773: out <= 16'h03E7;    16'd58774: out <= 16'h0375;    16'd58775: out <= 16'h09F9;
    16'd58776: out <= 16'h028D;    16'd58777: out <= 16'h018A;    16'd58778: out <= 16'h0413;    16'd58779: out <= 16'h0438;
    16'd58780: out <= 16'hFE56;    16'd58781: out <= 16'h0039;    16'd58782: out <= 16'hFF62;    16'd58783: out <= 16'h0233;
    16'd58784: out <= 16'h04B3;    16'd58785: out <= 16'h03C4;    16'd58786: out <= 16'h0440;    16'd58787: out <= 16'h095F;
    16'd58788: out <= 16'h04D2;    16'd58789: out <= 16'h02FD;    16'd58790: out <= 16'h077D;    16'd58791: out <= 16'hFEF9;
    16'd58792: out <= 16'h032F;    16'd58793: out <= 16'h0905;    16'd58794: out <= 16'hFFE4;    16'd58795: out <= 16'h0406;
    16'd58796: out <= 16'h039A;    16'd58797: out <= 16'h06CF;    16'd58798: out <= 16'h056E;    16'd58799: out <= 16'h061F;
    16'd58800: out <= 16'h023B;    16'd58801: out <= 16'hFFC1;    16'd58802: out <= 16'h042A;    16'd58803: out <= 16'h0280;
    16'd58804: out <= 16'h0519;    16'd58805: out <= 16'h0146;    16'd58806: out <= 16'h096E;    16'd58807: out <= 16'h02F4;
    16'd58808: out <= 16'h07A5;    16'd58809: out <= 16'h02E9;    16'd58810: out <= 16'h055A;    16'd58811: out <= 16'h0795;
    16'd58812: out <= 16'h06CD;    16'd58813: out <= 16'h044B;    16'd58814: out <= 16'h019C;    16'd58815: out <= 16'h094E;
    16'd58816: out <= 16'h0A60;    16'd58817: out <= 16'hFFD4;    16'd58818: out <= 16'h0681;    16'd58819: out <= 16'h0030;
    16'd58820: out <= 16'h03C9;    16'd58821: out <= 16'h083C;    16'd58822: out <= 16'h0581;    16'd58823: out <= 16'h01E4;
    16'd58824: out <= 16'h08EC;    16'd58825: out <= 16'h0001;    16'd58826: out <= 16'h02EE;    16'd58827: out <= 16'h03BD;
    16'd58828: out <= 16'h00C1;    16'd58829: out <= 16'hFFE8;    16'd58830: out <= 16'hFFBC;    16'd58831: out <= 16'hFF83;
    16'd58832: out <= 16'h013D;    16'd58833: out <= 16'hF705;    16'd58834: out <= 16'h03B8;    16'd58835: out <= 16'h027D;
    16'd58836: out <= 16'hF9B3;    16'd58837: out <= 16'hFBFE;    16'd58838: out <= 16'hFD85;    16'd58839: out <= 16'hFD5D;
    16'd58840: out <= 16'hFE4D;    16'd58841: out <= 16'hFBF5;    16'd58842: out <= 16'h0223;    16'd58843: out <= 16'h0187;
    16'd58844: out <= 16'hFF66;    16'd58845: out <= 16'hFECE;    16'd58846: out <= 16'hFFAB;    16'd58847: out <= 16'hFEE0;
    16'd58848: out <= 16'h034D;    16'd58849: out <= 16'hFCD3;    16'd58850: out <= 16'hFD79;    16'd58851: out <= 16'hFBDD;
    16'd58852: out <= 16'hFA46;    16'd58853: out <= 16'hFF66;    16'd58854: out <= 16'hFCC3;    16'd58855: out <= 16'h01DD;
    16'd58856: out <= 16'h0027;    16'd58857: out <= 16'hFBF1;    16'd58858: out <= 16'hFC48;    16'd58859: out <= 16'hFDF7;
    16'd58860: out <= 16'hFFF1;    16'd58861: out <= 16'h037E;    16'd58862: out <= 16'h081B;    16'd58863: out <= 16'h0100;
    16'd58864: out <= 16'h07B0;    16'd58865: out <= 16'hFB71;    16'd58866: out <= 16'hFA67;    16'd58867: out <= 16'hFB23;
    16'd58868: out <= 16'hFEA0;    16'd58869: out <= 16'h0055;    16'd58870: out <= 16'hFDE2;    16'd58871: out <= 16'h014C;
    16'd58872: out <= 16'h0147;    16'd58873: out <= 16'hFF2A;    16'd58874: out <= 16'h0497;    16'd58875: out <= 16'hFBD4;
    16'd58876: out <= 16'hFEEB;    16'd58877: out <= 16'hF912;    16'd58878: out <= 16'hF7B1;    16'd58879: out <= 16'h042F;
    16'd58880: out <= 16'h0044;    16'd58881: out <= 16'hFDF4;    16'd58882: out <= 16'h0145;    16'd58883: out <= 16'hFB06;
    16'd58884: out <= 16'h0225;    16'd58885: out <= 16'h0089;    16'd58886: out <= 16'h023D;    16'd58887: out <= 16'h0183;
    16'd58888: out <= 16'h06F8;    16'd58889: out <= 16'h03B2;    16'd58890: out <= 16'hFEE4;    16'd58891: out <= 16'h06C9;
    16'd58892: out <= 16'hFF8B;    16'd58893: out <= 16'h02E5;    16'd58894: out <= 16'h019E;    16'd58895: out <= 16'h06FC;
    16'd58896: out <= 16'hFB56;    16'd58897: out <= 16'h002A;    16'd58898: out <= 16'hFDB3;    16'd58899: out <= 16'h00AB;
    16'd58900: out <= 16'h0083;    16'd58901: out <= 16'hFCA5;    16'd58902: out <= 16'hFF63;    16'd58903: out <= 16'hFFE3;
    16'd58904: out <= 16'hFBD2;    16'd58905: out <= 16'hFF7F;    16'd58906: out <= 16'hFFE7;    16'd58907: out <= 16'hFA4E;
    16'd58908: out <= 16'hFE92;    16'd58909: out <= 16'h0166;    16'd58910: out <= 16'h0100;    16'd58911: out <= 16'h02AA;
    16'd58912: out <= 16'h028B;    16'd58913: out <= 16'h0110;    16'd58914: out <= 16'hFDA9;    16'd58915: out <= 16'hFDF4;
    16'd58916: out <= 16'h0126;    16'd58917: out <= 16'hFEBF;    16'd58918: out <= 16'hFE34;    16'd58919: out <= 16'h028F;
    16'd58920: out <= 16'hFB8C;    16'd58921: out <= 16'h00BD;    16'd58922: out <= 16'hFD04;    16'd58923: out <= 16'h013F;
    16'd58924: out <= 16'hFF91;    16'd58925: out <= 16'hFD7D;    16'd58926: out <= 16'h0553;    16'd58927: out <= 16'h043E;
    16'd58928: out <= 16'h036F;    16'd58929: out <= 16'h03C3;    16'd58930: out <= 16'h0435;    16'd58931: out <= 16'hFFED;
    16'd58932: out <= 16'h0820;    16'd58933: out <= 16'h031A;    16'd58934: out <= 16'h09E5;    16'd58935: out <= 16'h01AF;
    16'd58936: out <= 16'h0680;    16'd58937: out <= 16'hFBA5;    16'd58938: out <= 16'h087A;    16'd58939: out <= 16'h054D;
    16'd58940: out <= 16'h067F;    16'd58941: out <= 16'h06E0;    16'd58942: out <= 16'hFD6D;    16'd58943: out <= 16'h0259;
    16'd58944: out <= 16'h02E5;    16'd58945: out <= 16'h0076;    16'd58946: out <= 16'h0406;    16'd58947: out <= 16'h0332;
    16'd58948: out <= 16'h03B7;    16'd58949: out <= 16'h0D61;    16'd58950: out <= 16'h0505;    16'd58951: out <= 16'h0687;
    16'd58952: out <= 16'hFF19;    16'd58953: out <= 16'hFA7A;    16'd58954: out <= 16'h05B9;    16'd58955: out <= 16'h07EC;
    16'd58956: out <= 16'h0A44;    16'd58957: out <= 16'h01E2;    16'd58958: out <= 16'h037A;    16'd58959: out <= 16'h0536;
    16'd58960: out <= 16'h020B;    16'd58961: out <= 16'hFDF3;    16'd58962: out <= 16'hFFA3;    16'd58963: out <= 16'hFE6C;
    16'd58964: out <= 16'h04B9;    16'd58965: out <= 16'h018C;    16'd58966: out <= 16'hFC13;    16'd58967: out <= 16'h00EC;
    16'd58968: out <= 16'h048D;    16'd58969: out <= 16'h005D;    16'd58970: out <= 16'h05B3;    16'd58971: out <= 16'h08DD;
    16'd58972: out <= 16'h06F7;    16'd58973: out <= 16'hFE98;    16'd58974: out <= 16'h0050;    16'd58975: out <= 16'hFF57;
    16'd58976: out <= 16'h05E0;    16'd58977: out <= 16'h08CA;    16'd58978: out <= 16'h08C7;    16'd58979: out <= 16'h0E7C;
    16'd58980: out <= 16'h0697;    16'd58981: out <= 16'h0388;    16'd58982: out <= 16'h01D7;    16'd58983: out <= 16'h0365;
    16'd58984: out <= 16'hFD31;    16'd58985: out <= 16'hFE29;    16'd58986: out <= 16'h092C;    16'd58987: out <= 16'h04D7;
    16'd58988: out <= 16'h09D4;    16'd58989: out <= 16'h05DF;    16'd58990: out <= 16'h030B;    16'd58991: out <= 16'h07F7;
    16'd58992: out <= 16'h04EF;    16'd58993: out <= 16'h032F;    16'd58994: out <= 16'h0B73;    16'd58995: out <= 16'h0021;
    16'd58996: out <= 16'h02CB;    16'd58997: out <= 16'h0479;    16'd58998: out <= 16'h01EC;    16'd58999: out <= 16'h04B2;
    16'd59000: out <= 16'h03C9;    16'd59001: out <= 16'h02B6;    16'd59002: out <= 16'hFF77;    16'd59003: out <= 16'h02DC;
    16'd59004: out <= 16'h0693;    16'd59005: out <= 16'h01CB;    16'd59006: out <= 16'hFF87;    16'd59007: out <= 16'h066B;
    16'd59008: out <= 16'h0602;    16'd59009: out <= 16'hFEAF;    16'd59010: out <= 16'h0457;    16'd59011: out <= 16'h0AA1;
    16'd59012: out <= 16'h0543;    16'd59013: out <= 16'h03CC;    16'd59014: out <= 16'h015C;    16'd59015: out <= 16'h00E4;
    16'd59016: out <= 16'h00D6;    16'd59017: out <= 16'h045B;    16'd59018: out <= 16'h0BED;    16'd59019: out <= 16'hFF98;
    16'd59020: out <= 16'h0514;    16'd59021: out <= 16'h0854;    16'd59022: out <= 16'h00F1;    16'd59023: out <= 16'h037E;
    16'd59024: out <= 16'h04A9;    16'd59025: out <= 16'h03AB;    16'd59026: out <= 16'h0C02;    16'd59027: out <= 16'h0369;
    16'd59028: out <= 16'h01EF;    16'd59029: out <= 16'h04B4;    16'd59030: out <= 16'h04C9;    16'd59031: out <= 16'hFCDF;
    16'd59032: out <= 16'h058B;    16'd59033: out <= 16'h012D;    16'd59034: out <= 16'hFD1A;    16'd59035: out <= 16'h0492;
    16'd59036: out <= 16'h021A;    16'd59037: out <= 16'h00F7;    16'd59038: out <= 16'h0A8B;    16'd59039: out <= 16'h0512;
    16'd59040: out <= 16'h03FC;    16'd59041: out <= 16'h0877;    16'd59042: out <= 16'h089B;    16'd59043: out <= 16'h0BF1;
    16'd59044: out <= 16'h0374;    16'd59045: out <= 16'h0975;    16'd59046: out <= 16'h09C3;    16'd59047: out <= 16'h06B2;
    16'd59048: out <= 16'h0186;    16'd59049: out <= 16'h01F8;    16'd59050: out <= 16'h0001;    16'd59051: out <= 16'hFF09;
    16'd59052: out <= 16'h03CF;    16'd59053: out <= 16'hFFE6;    16'd59054: out <= 16'hFD9C;    16'd59055: out <= 16'h0190;
    16'd59056: out <= 16'h0A65;    16'd59057: out <= 16'h082C;    16'd59058: out <= 16'hFD1E;    16'd59059: out <= 16'h044A;
    16'd59060: out <= 16'h0AA5;    16'd59061: out <= 16'h0588;    16'd59062: out <= 16'h0198;    16'd59063: out <= 16'h04F1;
    16'd59064: out <= 16'h04A8;    16'd59065: out <= 16'hFFA1;    16'd59066: out <= 16'h0620;    16'd59067: out <= 16'h01E2;
    16'd59068: out <= 16'h03BB;    16'd59069: out <= 16'h0752;    16'd59070: out <= 16'h0770;    16'd59071: out <= 16'h013C;
    16'd59072: out <= 16'h0668;    16'd59073: out <= 16'h01AE;    16'd59074: out <= 16'h0309;    16'd59075: out <= 16'h008F;
    16'd59076: out <= 16'h00E7;    16'd59077: out <= 16'h0263;    16'd59078: out <= 16'h0021;    16'd59079: out <= 16'h00DC;
    16'd59080: out <= 16'hFDE0;    16'd59081: out <= 16'hFA19;    16'd59082: out <= 16'h02FF;    16'd59083: out <= 16'hFE28;
    16'd59084: out <= 16'h027A;    16'd59085: out <= 16'h0345;    16'd59086: out <= 16'hFD32;    16'd59087: out <= 16'hFC77;
    16'd59088: out <= 16'h00BA;    16'd59089: out <= 16'hFBA9;    16'd59090: out <= 16'hFD58;    16'd59091: out <= 16'h029C;
    16'd59092: out <= 16'hF895;    16'd59093: out <= 16'h02E4;    16'd59094: out <= 16'hFF54;    16'd59095: out <= 16'h008C;
    16'd59096: out <= 16'h0019;    16'd59097: out <= 16'h0719;    16'd59098: out <= 16'hFE36;    16'd59099: out <= 16'hFD04;
    16'd59100: out <= 16'hFE8E;    16'd59101: out <= 16'h0A9C;    16'd59102: out <= 16'hFEA4;    16'd59103: out <= 16'hFC9B;
    16'd59104: out <= 16'h015A;    16'd59105: out <= 16'hFEF3;    16'd59106: out <= 16'hFF6F;    16'd59107: out <= 16'h0570;
    16'd59108: out <= 16'hFE83;    16'd59109: out <= 16'hFBC3;    16'd59110: out <= 16'h025E;    16'd59111: out <= 16'hFF45;
    16'd59112: out <= 16'h0416;    16'd59113: out <= 16'hFE49;    16'd59114: out <= 16'h0266;    16'd59115: out <= 16'hFF34;
    16'd59116: out <= 16'hFD83;    16'd59117: out <= 16'hFBF1;    16'd59118: out <= 16'h030D;    16'd59119: out <= 16'hFC0E;
    16'd59120: out <= 16'hFF83;    16'd59121: out <= 16'h081A;    16'd59122: out <= 16'hF8AB;    16'd59123: out <= 16'hFCA1;
    16'd59124: out <= 16'hFCA5;    16'd59125: out <= 16'hFF95;    16'd59126: out <= 16'hFBAE;    16'd59127: out <= 16'hFBAA;
    16'd59128: out <= 16'hF69D;    16'd59129: out <= 16'hFBFF;    16'd59130: out <= 16'h0804;    16'd59131: out <= 16'h0046;
    16'd59132: out <= 16'h0106;    16'd59133: out <= 16'h00C5;    16'd59134: out <= 16'hF90D;    16'd59135: out <= 16'h0165;
    16'd59136: out <= 16'h00BC;    16'd59137: out <= 16'hFE9C;    16'd59138: out <= 16'hFFC6;    16'd59139: out <= 16'hFD57;
    16'd59140: out <= 16'hFFE3;    16'd59141: out <= 16'h006B;    16'd59142: out <= 16'h0287;    16'd59143: out <= 16'h0158;
    16'd59144: out <= 16'h0303;    16'd59145: out <= 16'h01D9;    16'd59146: out <= 16'h076B;    16'd59147: out <= 16'h02E6;
    16'd59148: out <= 16'h00D2;    16'd59149: out <= 16'hFF51;    16'd59150: out <= 16'hF8D9;    16'd59151: out <= 16'hFBE6;
    16'd59152: out <= 16'h050E;    16'd59153: out <= 16'h0032;    16'd59154: out <= 16'h0181;    16'd59155: out <= 16'h047F;
    16'd59156: out <= 16'h060B;    16'd59157: out <= 16'h00C2;    16'd59158: out <= 16'h02A1;    16'd59159: out <= 16'h044F;
    16'd59160: out <= 16'hFDFD;    16'd59161: out <= 16'hFFD6;    16'd59162: out <= 16'h004C;    16'd59163: out <= 16'h0512;
    16'd59164: out <= 16'h03AD;    16'd59165: out <= 16'hFD32;    16'd59166: out <= 16'hFCE8;    16'd59167: out <= 16'h0236;
    16'd59168: out <= 16'h00EC;    16'd59169: out <= 16'hFCAF;    16'd59170: out <= 16'hFDA8;    16'd59171: out <= 16'h02F4;
    16'd59172: out <= 16'hFF01;    16'd59173: out <= 16'h038B;    16'd59174: out <= 16'hFFF5;    16'd59175: out <= 16'hFDD8;
    16'd59176: out <= 16'h01F1;    16'd59177: out <= 16'hFB1C;    16'd59178: out <= 16'hFAF7;    16'd59179: out <= 16'hFFFD;
    16'd59180: out <= 16'h02A9;    16'd59181: out <= 16'h010D;    16'd59182: out <= 16'hFA13;    16'd59183: out <= 16'h02F5;
    16'd59184: out <= 16'h03D8;    16'd59185: out <= 16'h0008;    16'd59186: out <= 16'h0E20;    16'd59187: out <= 16'h0723;
    16'd59188: out <= 16'h0849;    16'd59189: out <= 16'h09DD;    16'd59190: out <= 16'h057E;    16'd59191: out <= 16'h07E0;
    16'd59192: out <= 16'h0852;    16'd59193: out <= 16'h003A;    16'd59194: out <= 16'h010D;    16'd59195: out <= 16'h006F;
    16'd59196: out <= 16'h03CA;    16'd59197: out <= 16'h0747;    16'd59198: out <= 16'h043D;    16'd59199: out <= 16'h0008;
    16'd59200: out <= 16'hFFBE;    16'd59201: out <= 16'h0679;    16'd59202: out <= 16'h03DF;    16'd59203: out <= 16'h0427;
    16'd59204: out <= 16'h02EB;    16'd59205: out <= 16'h0378;    16'd59206: out <= 16'h0793;    16'd59207: out <= 16'h0880;
    16'd59208: out <= 16'h00ED;    16'd59209: out <= 16'h08E4;    16'd59210: out <= 16'h0B09;    16'd59211: out <= 16'h068A;
    16'd59212: out <= 16'h027D;    16'd59213: out <= 16'h06E4;    16'd59214: out <= 16'h03E8;    16'd59215: out <= 16'h050D;
    16'd59216: out <= 16'h078D;    16'd59217: out <= 16'h0178;    16'd59218: out <= 16'h05BD;    16'd59219: out <= 16'h01D6;
    16'd59220: out <= 16'hFBA3;    16'd59221: out <= 16'h03B4;    16'd59222: out <= 16'h01FA;    16'd59223: out <= 16'h03B6;
    16'd59224: out <= 16'h02C2;    16'd59225: out <= 16'h036D;    16'd59226: out <= 16'h03A3;    16'd59227: out <= 16'hFEB5;
    16'd59228: out <= 16'h0984;    16'd59229: out <= 16'h0390;    16'd59230: out <= 16'h047E;    16'd59231: out <= 16'h019C;
    16'd59232: out <= 16'h040C;    16'd59233: out <= 16'h0350;    16'd59234: out <= 16'h0758;    16'd59235: out <= 16'h03E2;
    16'd59236: out <= 16'h058E;    16'd59237: out <= 16'hFEFA;    16'd59238: out <= 16'h002F;    16'd59239: out <= 16'h06E0;
    16'd59240: out <= 16'h021F;    16'd59241: out <= 16'h02A1;    16'd59242: out <= 16'h050A;    16'd59243: out <= 16'hFC3C;
    16'd59244: out <= 16'h012C;    16'd59245: out <= 16'h01DF;    16'd59246: out <= 16'h01F9;    16'd59247: out <= 16'h0439;
    16'd59248: out <= 16'h024D;    16'd59249: out <= 16'h02FC;    16'd59250: out <= 16'h01DE;    16'd59251: out <= 16'h074E;
    16'd59252: out <= 16'hFBE3;    16'd59253: out <= 16'h025C;    16'd59254: out <= 16'h063A;    16'd59255: out <= 16'h052C;
    16'd59256: out <= 16'h0268;    16'd59257: out <= 16'h096A;    16'd59258: out <= 16'h0229;    16'd59259: out <= 16'h0158;
    16'd59260: out <= 16'h0735;    16'd59261: out <= 16'h021B;    16'd59262: out <= 16'h0188;    16'd59263: out <= 16'h0536;
    16'd59264: out <= 16'h0856;    16'd59265: out <= 16'h06AF;    16'd59266: out <= 16'h0433;    16'd59267: out <= 16'hFDB8;
    16'd59268: out <= 16'h03B4;    16'd59269: out <= 16'hFE0B;    16'd59270: out <= 16'h05C5;    16'd59271: out <= 16'h00B6;
    16'd59272: out <= 16'h058C;    16'd59273: out <= 16'h0014;    16'd59274: out <= 16'h03BA;    16'd59275: out <= 16'h07A1;
    16'd59276: out <= 16'h03D6;    16'd59277: out <= 16'h07F0;    16'd59278: out <= 16'h099F;    16'd59279: out <= 16'h06AC;
    16'd59280: out <= 16'h02BC;    16'd59281: out <= 16'hFDC3;    16'd59282: out <= 16'hFF17;    16'd59283: out <= 16'h0752;
    16'd59284: out <= 16'h0296;    16'd59285: out <= 16'h0475;    16'd59286: out <= 16'hFE7A;    16'd59287: out <= 16'h088F;
    16'd59288: out <= 16'h0514;    16'd59289: out <= 16'h0277;    16'd59290: out <= 16'h0832;    16'd59291: out <= 16'h043C;
    16'd59292: out <= 16'hFD4B;    16'd59293: out <= 16'h0493;    16'd59294: out <= 16'h0228;    16'd59295: out <= 16'h0565;
    16'd59296: out <= 16'h0520;    16'd59297: out <= 16'h05E2;    16'd59298: out <= 16'h0BCF;    16'd59299: out <= 16'h072F;
    16'd59300: out <= 16'h003E;    16'd59301: out <= 16'h02DE;    16'd59302: out <= 16'h0522;    16'd59303: out <= 16'h0350;
    16'd59304: out <= 16'hFFA6;    16'd59305: out <= 16'h0613;    16'd59306: out <= 16'hFC3F;    16'd59307: out <= 16'h0432;
    16'd59308: out <= 16'h0182;    16'd59309: out <= 16'h030F;    16'd59310: out <= 16'h0569;    16'd59311: out <= 16'hFCAE;
    16'd59312: out <= 16'hFF59;    16'd59313: out <= 16'hFA8E;    16'd59314: out <= 16'h0119;    16'd59315: out <= 16'h0738;
    16'd59316: out <= 16'h05F1;    16'd59317: out <= 16'h04F7;    16'd59318: out <= 16'h0709;    16'd59319: out <= 16'h015C;
    16'd59320: out <= 16'h04C4;    16'd59321: out <= 16'hFD3C;    16'd59322: out <= 16'h0378;    16'd59323: out <= 16'hFC8D;
    16'd59324: out <= 16'h0437;    16'd59325: out <= 16'h0586;    16'd59326: out <= 16'h0330;    16'd59327: out <= 16'h09C2;
    16'd59328: out <= 16'h04CC;    16'd59329: out <= 16'h08B0;    16'd59330: out <= 16'h0216;    16'd59331: out <= 16'hFBC3;
    16'd59332: out <= 16'hFC97;    16'd59333: out <= 16'h0773;    16'd59334: out <= 16'h0429;    16'd59335: out <= 16'hFEB5;
    16'd59336: out <= 16'hFEEA;    16'd59337: out <= 16'h00D8;    16'd59338: out <= 16'hFC0F;    16'd59339: out <= 16'h05F9;
    16'd59340: out <= 16'hFEDC;    16'd59341: out <= 16'hFF4E;    16'd59342: out <= 16'h0163;    16'd59343: out <= 16'h01D5;
    16'd59344: out <= 16'hFF8F;    16'd59345: out <= 16'h02FE;    16'd59346: out <= 16'h0433;    16'd59347: out <= 16'hFA85;
    16'd59348: out <= 16'h04FA;    16'd59349: out <= 16'hF9E4;    16'd59350: out <= 16'h0041;    16'd59351: out <= 16'h046C;
    16'd59352: out <= 16'hFA6F;    16'd59353: out <= 16'h0159;    16'd59354: out <= 16'h0372;    16'd59355: out <= 16'hFF7F;
    16'd59356: out <= 16'h004B;    16'd59357: out <= 16'h04A2;    16'd59358: out <= 16'h0018;    16'd59359: out <= 16'h0081;
    16'd59360: out <= 16'hFDE8;    16'd59361: out <= 16'hF784;    16'd59362: out <= 16'h054F;    16'd59363: out <= 16'hFD32;
    16'd59364: out <= 16'h0077;    16'd59365: out <= 16'hF9B1;    16'd59366: out <= 16'h004E;    16'd59367: out <= 16'hFFC2;
    16'd59368: out <= 16'hFDB7;    16'd59369: out <= 16'hFDA7;    16'd59370: out <= 16'h0090;    16'd59371: out <= 16'h02D3;
    16'd59372: out <= 16'h028C;    16'd59373: out <= 16'h04A8;    16'd59374: out <= 16'h0714;    16'd59375: out <= 16'h0305;
    16'd59376: out <= 16'hFD89;    16'd59377: out <= 16'h01F3;    16'd59378: out <= 16'h0652;    16'd59379: out <= 16'h006E;
    16'd59380: out <= 16'hFE4A;    16'd59381: out <= 16'hFB08;    16'd59382: out <= 16'h02F8;    16'd59383: out <= 16'h0044;
    16'd59384: out <= 16'h01AC;    16'd59385: out <= 16'h035B;    16'd59386: out <= 16'h0717;    16'd59387: out <= 16'h022F;
    16'd59388: out <= 16'hFCDA;    16'd59389: out <= 16'h06D4;    16'd59390: out <= 16'h0411;    16'd59391: out <= 16'h0035;
    16'd59392: out <= 16'hFBCE;    16'd59393: out <= 16'hFDED;    16'd59394: out <= 16'hFE78;    16'd59395: out <= 16'h02CA;
    16'd59396: out <= 16'h04C3;    16'd59397: out <= 16'hFC2E;    16'd59398: out <= 16'hFE11;    16'd59399: out <= 16'hFBE3;
    16'd59400: out <= 16'hFF46;    16'd59401: out <= 16'hFFF2;    16'd59402: out <= 16'hFDD9;    16'd59403: out <= 16'hFDB0;
    16'd59404: out <= 16'h0098;    16'd59405: out <= 16'hFBB5;    16'd59406: out <= 16'h01FE;    16'd59407: out <= 16'hFFBE;
    16'd59408: out <= 16'hFFD7;    16'd59409: out <= 16'h024F;    16'd59410: out <= 16'h0341;    16'd59411: out <= 16'h01F4;
    16'd59412: out <= 16'hFF1D;    16'd59413: out <= 16'hFE9F;    16'd59414: out <= 16'hFF65;    16'd59415: out <= 16'hF6C4;
    16'd59416: out <= 16'h016A;    16'd59417: out <= 16'h0680;    16'd59418: out <= 16'h0452;    16'd59419: out <= 16'hFD24;
    16'd59420: out <= 16'hFEA2;    16'd59421: out <= 16'hFD29;    16'd59422: out <= 16'hFB49;    16'd59423: out <= 16'h0586;
    16'd59424: out <= 16'hFE2B;    16'd59425: out <= 16'h00C1;    16'd59426: out <= 16'hF8D1;    16'd59427: out <= 16'hFC80;
    16'd59428: out <= 16'h0059;    16'd59429: out <= 16'hFA10;    16'd59430: out <= 16'h0211;    16'd59431: out <= 16'hFE4A;
    16'd59432: out <= 16'h05CC;    16'd59433: out <= 16'hFF80;    16'd59434: out <= 16'h01E0;    16'd59435: out <= 16'h0058;
    16'd59436: out <= 16'h029B;    16'd59437: out <= 16'h01A2;    16'd59438: out <= 16'hFE86;    16'd59439: out <= 16'h0414;
    16'd59440: out <= 16'h04EB;    16'd59441: out <= 16'h01DF;    16'd59442: out <= 16'h0587;    16'd59443: out <= 16'hFC27;
    16'd59444: out <= 16'h0B4E;    16'd59445: out <= 16'h0552;    16'd59446: out <= 16'h06C5;    16'd59447: out <= 16'h0083;
    16'd59448: out <= 16'h0256;    16'd59449: out <= 16'h01BD;    16'd59450: out <= 16'hFCD8;    16'd59451: out <= 16'h091D;
    16'd59452: out <= 16'h07C8;    16'd59453: out <= 16'hFF0D;    16'd59454: out <= 16'h05FF;    16'd59455: out <= 16'h0384;
    16'd59456: out <= 16'h0260;    16'd59457: out <= 16'h06A0;    16'd59458: out <= 16'h0379;    16'd59459: out <= 16'h0259;
    16'd59460: out <= 16'h03FC;    16'd59461: out <= 16'h0EE0;    16'd59462: out <= 16'h0877;    16'd59463: out <= 16'hFF39;
    16'd59464: out <= 16'h0939;    16'd59465: out <= 16'h009B;    16'd59466: out <= 16'hFDC2;    16'd59467: out <= 16'h0388;
    16'd59468: out <= 16'h0362;    16'd59469: out <= 16'hFC9A;    16'd59470: out <= 16'h0726;    16'd59471: out <= 16'h070A;
    16'd59472: out <= 16'h02BB;    16'd59473: out <= 16'h0C6B;    16'd59474: out <= 16'h112E;    16'd59475: out <= 16'h029A;
    16'd59476: out <= 16'h062D;    16'd59477: out <= 16'h0C32;    16'd59478: out <= 16'h0416;    16'd59479: out <= 16'h071C;
    16'd59480: out <= 16'h0250;    16'd59481: out <= 16'h0486;    16'd59482: out <= 16'h03C1;    16'd59483: out <= 16'h07C9;
    16'd59484: out <= 16'h04EC;    16'd59485: out <= 16'hFFED;    16'd59486: out <= 16'h024D;    16'd59487: out <= 16'hFFE6;
    16'd59488: out <= 16'h0A10;    16'd59489: out <= 16'h050D;    16'd59490: out <= 16'hFDAA;    16'd59491: out <= 16'h07BF;
    16'd59492: out <= 16'h067F;    16'd59493: out <= 16'hFEC8;    16'd59494: out <= 16'h0558;    16'd59495: out <= 16'h07A9;
    16'd59496: out <= 16'hF9E9;    16'd59497: out <= 16'hFD1C;    16'd59498: out <= 16'h01CE;    16'd59499: out <= 16'h002C;
    16'd59500: out <= 16'h030B;    16'd59501: out <= 16'h0180;    16'd59502: out <= 16'h027A;    16'd59503: out <= 16'h027C;
    16'd59504: out <= 16'h025D;    16'd59505: out <= 16'h0190;    16'd59506: out <= 16'h0766;    16'd59507: out <= 16'hFC1E;
    16'd59508: out <= 16'hFE7C;    16'd59509: out <= 16'hFFFA;    16'd59510: out <= 16'h0460;    16'd59511: out <= 16'h0B83;
    16'd59512: out <= 16'hFA2A;    16'd59513: out <= 16'h0152;    16'd59514: out <= 16'h06F7;    16'd59515: out <= 16'h02A6;
    16'd59516: out <= 16'h01CA;    16'd59517: out <= 16'hFF84;    16'd59518: out <= 16'h05A0;    16'd59519: out <= 16'h0286;
    16'd59520: out <= 16'hFFD6;    16'd59521: out <= 16'h07F3;    16'd59522: out <= 16'h02FD;    16'd59523: out <= 16'h0614;
    16'd59524: out <= 16'h0453;    16'd59525: out <= 16'h0596;    16'd59526: out <= 16'h05B1;    16'd59527: out <= 16'h02ED;
    16'd59528: out <= 16'h0592;    16'd59529: out <= 16'hFF47;    16'd59530: out <= 16'h012A;    16'd59531: out <= 16'h0796;
    16'd59532: out <= 16'h0A21;    16'd59533: out <= 16'h0380;    16'd59534: out <= 16'h09A9;    16'd59535: out <= 16'h05E3;
    16'd59536: out <= 16'h01A1;    16'd59537: out <= 16'hFFD9;    16'd59538: out <= 16'h0A3B;    16'd59539: out <= 16'h0882;
    16'd59540: out <= 16'h0A3D;    16'd59541: out <= 16'h0460;    16'd59542: out <= 16'h084A;    16'd59543: out <= 16'h0485;
    16'd59544: out <= 16'h041A;    16'd59545: out <= 16'h02E8;    16'd59546: out <= 16'h0500;    16'd59547: out <= 16'h020A;
    16'd59548: out <= 16'h041F;    16'd59549: out <= 16'h0698;    16'd59550: out <= 16'h06BA;    16'd59551: out <= 16'h0039;
    16'd59552: out <= 16'h0CC4;    16'd59553: out <= 16'h038C;    16'd59554: out <= 16'h068A;    16'd59555: out <= 16'hFF1A;
    16'd59556: out <= 16'hFE93;    16'd59557: out <= 16'h0A1F;    16'd59558: out <= 16'h05D5;    16'd59559: out <= 16'h06DE;
    16'd59560: out <= 16'h019B;    16'd59561: out <= 16'h0810;    16'd59562: out <= 16'h0060;    16'd59563: out <= 16'h0195;
    16'd59564: out <= 16'h036F;    16'd59565: out <= 16'hFC83;    16'd59566: out <= 16'h0636;    16'd59567: out <= 16'h089F;
    16'd59568: out <= 16'h037B;    16'd59569: out <= 16'h0426;    16'd59570: out <= 16'hFEE9;    16'd59571: out <= 16'h050F;
    16'd59572: out <= 16'h0782;    16'd59573: out <= 16'hFF85;    16'd59574: out <= 16'h000D;    16'd59575: out <= 16'h08C4;
    16'd59576: out <= 16'h041C;    16'd59577: out <= 16'hFA8F;    16'd59578: out <= 16'h0E28;    16'd59579: out <= 16'h0619;
    16'd59580: out <= 16'h0161;    16'd59581: out <= 16'h057A;    16'd59582: out <= 16'hFF79;    16'd59583: out <= 16'hFFBA;
    16'd59584: out <= 16'h055E;    16'd59585: out <= 16'h0460;    16'd59586: out <= 16'h05AA;    16'd59587: out <= 16'h000D;
    16'd59588: out <= 16'h00D0;    16'd59589: out <= 16'h04C9;    16'd59590: out <= 16'h06C0;    16'd59591: out <= 16'h01FD;
    16'd59592: out <= 16'h02F6;    16'd59593: out <= 16'h0516;    16'd59594: out <= 16'h085B;    16'd59595: out <= 16'h0474;
    16'd59596: out <= 16'h04BD;    16'd59597: out <= 16'hFDD2;    16'd59598: out <= 16'h00C8;    16'd59599: out <= 16'h0115;
    16'd59600: out <= 16'hF902;    16'd59601: out <= 16'hFC53;    16'd59602: out <= 16'hF8A4;    16'd59603: out <= 16'hF9FB;
    16'd59604: out <= 16'hFD10;    16'd59605: out <= 16'hFD00;    16'd59606: out <= 16'h00E7;    16'd59607: out <= 16'hF839;
    16'd59608: out <= 16'h008E;    16'd59609: out <= 16'h03D4;    16'd59610: out <= 16'h0115;    16'd59611: out <= 16'h012B;
    16'd59612: out <= 16'h00E2;    16'd59613: out <= 16'h01D8;    16'd59614: out <= 16'hFF21;    16'd59615: out <= 16'hFB52;
    16'd59616: out <= 16'h04E5;    16'd59617: out <= 16'hFDC3;    16'd59618: out <= 16'h05F5;    16'd59619: out <= 16'hF8A5;
    16'd59620: out <= 16'h01E1;    16'd59621: out <= 16'hFE29;    16'd59622: out <= 16'h0069;    16'd59623: out <= 16'h0162;
    16'd59624: out <= 16'h02DD;    16'd59625: out <= 16'hFBE7;    16'd59626: out <= 16'h0291;    16'd59627: out <= 16'h064B;
    16'd59628: out <= 16'hFF0A;    16'd59629: out <= 16'hF684;    16'd59630: out <= 16'h0297;    16'd59631: out <= 16'hFAA9;
    16'd59632: out <= 16'hFA94;    16'd59633: out <= 16'hFEB0;    16'd59634: out <= 16'h035D;    16'd59635: out <= 16'h0435;
    16'd59636: out <= 16'h061A;    16'd59637: out <= 16'h01F4;    16'd59638: out <= 16'hF9E1;    16'd59639: out <= 16'hFD15;
    16'd59640: out <= 16'h035E;    16'd59641: out <= 16'h005F;    16'd59642: out <= 16'hFED6;    16'd59643: out <= 16'hFAF0;
    16'd59644: out <= 16'hFEF5;    16'd59645: out <= 16'h0625;    16'd59646: out <= 16'h017A;    16'd59647: out <= 16'hFC24;
    16'd59648: out <= 16'h016D;    16'd59649: out <= 16'h0369;    16'd59650: out <= 16'h0202;    16'd59651: out <= 16'hFBBB;
    16'd59652: out <= 16'hFEAF;    16'd59653: out <= 16'h02C8;    16'd59654: out <= 16'h03B5;    16'd59655: out <= 16'h0628;
    16'd59656: out <= 16'h0185;    16'd59657: out <= 16'hFF8B;    16'd59658: out <= 16'hF9A3;    16'd59659: out <= 16'h043A;
    16'd59660: out <= 16'hF71D;    16'd59661: out <= 16'h0169;    16'd59662: out <= 16'h067D;    16'd59663: out <= 16'hFFD2;
    16'd59664: out <= 16'h02AB;    16'd59665: out <= 16'h007D;    16'd59666: out <= 16'hF9E4;    16'd59667: out <= 16'h05E9;
    16'd59668: out <= 16'h01B9;    16'd59669: out <= 16'h0181;    16'd59670: out <= 16'h0195;    16'd59671: out <= 16'h00DA;
    16'd59672: out <= 16'hFB59;    16'd59673: out <= 16'h0648;    16'd59674: out <= 16'h05D6;    16'd59675: out <= 16'h0099;
    16'd59676: out <= 16'hFBFE;    16'd59677: out <= 16'h0218;    16'd59678: out <= 16'hFC35;    16'd59679: out <= 16'h0076;
    16'd59680: out <= 16'hFB02;    16'd59681: out <= 16'hFB0F;    16'd59682: out <= 16'hFC72;    16'd59683: out <= 16'h00DD;
    16'd59684: out <= 16'hFB6A;    16'd59685: out <= 16'hF784;    16'd59686: out <= 16'hF880;    16'd59687: out <= 16'h0459;
    16'd59688: out <= 16'hFD21;    16'd59689: out <= 16'hFD86;    16'd59690: out <= 16'h07FA;    16'd59691: out <= 16'h027D;
    16'd59692: out <= 16'h0658;    16'd59693: out <= 16'hF8C1;    16'd59694: out <= 16'h0583;    16'd59695: out <= 16'h0206;
    16'd59696: out <= 16'h020C;    16'd59697: out <= 16'h00D4;    16'd59698: out <= 16'h0564;    16'd59699: out <= 16'h032B;
    16'd59700: out <= 16'h0404;    16'd59701: out <= 16'hFF6A;    16'd59702: out <= 16'h00A1;    16'd59703: out <= 16'h01B3;
    16'd59704: out <= 16'h0194;    16'd59705: out <= 16'hFFD2;    16'd59706: out <= 16'h055D;    16'd59707: out <= 16'h059C;
    16'd59708: out <= 16'h0756;    16'd59709: out <= 16'h05D6;    16'd59710: out <= 16'h05A3;    16'd59711: out <= 16'h01A4;
    16'd59712: out <= 16'h0013;    16'd59713: out <= 16'h053B;    16'd59714: out <= 16'h00D3;    16'd59715: out <= 16'h04DE;
    16'd59716: out <= 16'h04F5;    16'd59717: out <= 16'h0305;    16'd59718: out <= 16'h0938;    16'd59719: out <= 16'h012D;
    16'd59720: out <= 16'h0732;    16'd59721: out <= 16'h075A;    16'd59722: out <= 16'h0620;    16'd59723: out <= 16'h0641;
    16'd59724: out <= 16'hFF31;    16'd59725: out <= 16'h0289;    16'd59726: out <= 16'h00CA;    16'd59727: out <= 16'h03C7;
    16'd59728: out <= 16'h08B3;    16'd59729: out <= 16'h05B5;    16'd59730: out <= 16'h09DB;    16'd59731: out <= 16'h034D;
    16'd59732: out <= 16'h0669;    16'd59733: out <= 16'h0069;    16'd59734: out <= 16'h028E;    16'd59735: out <= 16'h00B7;
    16'd59736: out <= 16'h050D;    16'd59737: out <= 16'h0511;    16'd59738: out <= 16'hFD30;    16'd59739: out <= 16'h03F6;
    16'd59740: out <= 16'h02AC;    16'd59741: out <= 16'h045E;    16'd59742: out <= 16'hFFDD;    16'd59743: out <= 16'h0311;
    16'd59744: out <= 16'hFC02;    16'd59745: out <= 16'h06BD;    16'd59746: out <= 16'h03CA;    16'd59747: out <= 16'hF64F;
    16'd59748: out <= 16'hF76E;    16'd59749: out <= 16'h04A4;    16'd59750: out <= 16'hFED7;    16'd59751: out <= 16'h0251;
    16'd59752: out <= 16'hFDB5;    16'd59753: out <= 16'h04F6;    16'd59754: out <= 16'h00D5;    16'd59755: out <= 16'h077A;
    16'd59756: out <= 16'h0731;    16'd59757: out <= 16'hFE73;    16'd59758: out <= 16'hFDE4;    16'd59759: out <= 16'h039E;
    16'd59760: out <= 16'hFF8B;    16'd59761: out <= 16'hFE57;    16'd59762: out <= 16'hF96C;    16'd59763: out <= 16'h0029;
    16'd59764: out <= 16'h00F8;    16'd59765: out <= 16'h14AE;    16'd59766: out <= 16'h07F3;    16'd59767: out <= 16'h09B1;
    16'd59768: out <= 16'h017C;    16'd59769: out <= 16'h02D4;    16'd59770: out <= 16'hFE0B;    16'd59771: out <= 16'h074E;
    16'd59772: out <= 16'h033A;    16'd59773: out <= 16'h0083;    16'd59774: out <= 16'h01AB;    16'd59775: out <= 16'h060C;
    16'd59776: out <= 16'h0B83;    16'd59777: out <= 16'h06CF;    16'd59778: out <= 16'h067F;    16'd59779: out <= 16'h021C;
    16'd59780: out <= 16'h026D;    16'd59781: out <= 16'h0096;    16'd59782: out <= 16'h084F;    16'd59783: out <= 16'hFE76;
    16'd59784: out <= 16'h085B;    16'd59785: out <= 16'hFE9B;    16'd59786: out <= 16'h06F9;    16'd59787: out <= 16'h02E6;
    16'd59788: out <= 16'h08CB;    16'd59789: out <= 16'h0896;    16'd59790: out <= 16'h0195;    16'd59791: out <= 16'h090D;
    16'd59792: out <= 16'h04FF;    16'd59793: out <= 16'h0F72;    16'd59794: out <= 16'h03CE;    16'd59795: out <= 16'h0618;
    16'd59796: out <= 16'h02AA;    16'd59797: out <= 16'h0805;    16'd59798: out <= 16'h0AAB;    16'd59799: out <= 16'h0791;
    16'd59800: out <= 16'h035A;    16'd59801: out <= 16'h047C;    16'd59802: out <= 16'h0203;    16'd59803: out <= 16'h024E;
    16'd59804: out <= 16'h046C;    16'd59805: out <= 16'h0864;    16'd59806: out <= 16'hFA2E;    16'd59807: out <= 16'h0770;
    16'd59808: out <= 16'h01BE;    16'd59809: out <= 16'hFF49;    16'd59810: out <= 16'h07E8;    16'd59811: out <= 16'h07C9;
    16'd59812: out <= 16'h0D6C;    16'd59813: out <= 16'h05F7;    16'd59814: out <= 16'h097E;    16'd59815: out <= 16'h06AF;
    16'd59816: out <= 16'h04EF;    16'd59817: out <= 16'h00C0;    16'd59818: out <= 16'h0378;    16'd59819: out <= 16'h0918;
    16'd59820: out <= 16'h0267;    16'd59821: out <= 16'hFC0A;    16'd59822: out <= 16'h04D1;    16'd59823: out <= 16'hFF58;
    16'd59824: out <= 16'h05C2;    16'd59825: out <= 16'h05BF;    16'd59826: out <= 16'h021D;    16'd59827: out <= 16'hFD39;
    16'd59828: out <= 16'h01A0;    16'd59829: out <= 16'h0B37;    16'd59830: out <= 16'hF702;    16'd59831: out <= 16'hFDC1;
    16'd59832: out <= 16'h0545;    16'd59833: out <= 16'h04AA;    16'd59834: out <= 16'h0617;    16'd59835: out <= 16'h00FC;
    16'd59836: out <= 16'h0B28;    16'd59837: out <= 16'h0658;    16'd59838: out <= 16'h0136;    16'd59839: out <= 16'hFE2C;
    16'd59840: out <= 16'h0C70;    16'd59841: out <= 16'h026D;    16'd59842: out <= 16'h0573;    16'd59843: out <= 16'hFA8A;
    16'd59844: out <= 16'h02A6;    16'd59845: out <= 16'h0631;    16'd59846: out <= 16'hFE2C;    16'd59847: out <= 16'hFFEE;
    16'd59848: out <= 16'h01DD;    16'd59849: out <= 16'hF952;    16'd59850: out <= 16'hF98C;    16'd59851: out <= 16'hFC0A;
    16'd59852: out <= 16'h0779;    16'd59853: out <= 16'hFF8E;    16'd59854: out <= 16'h07FA;    16'd59855: out <= 16'h0573;
    16'd59856: out <= 16'h0697;    16'd59857: out <= 16'hFD1F;    16'd59858: out <= 16'h0315;    16'd59859: out <= 16'hFFC1;
    16'd59860: out <= 16'h0348;    16'd59861: out <= 16'hFDF7;    16'd59862: out <= 16'hFFEF;    16'd59863: out <= 16'h037C;
    16'd59864: out <= 16'h0749;    16'd59865: out <= 16'h01E8;    16'd59866: out <= 16'h058D;    16'd59867: out <= 16'hFBFA;
    16'd59868: out <= 16'h02B2;    16'd59869: out <= 16'hFC6D;    16'd59870: out <= 16'hFD1F;    16'd59871: out <= 16'h037C;
    16'd59872: out <= 16'h0340;    16'd59873: out <= 16'h04DF;    16'd59874: out <= 16'hFEC9;    16'd59875: out <= 16'hFE49;
    16'd59876: out <= 16'h015F;    16'd59877: out <= 16'h01C0;    16'd59878: out <= 16'h02D6;    16'd59879: out <= 16'h01A0;
    16'd59880: out <= 16'h000B;    16'd59881: out <= 16'h014F;    16'd59882: out <= 16'h01C9;    16'd59883: out <= 16'hFE02;
    16'd59884: out <= 16'hFA6D;    16'd59885: out <= 16'h0353;    16'd59886: out <= 16'h00D8;    16'd59887: out <= 16'h00B6;
    16'd59888: out <= 16'h0097;    16'd59889: out <= 16'hF901;    16'd59890: out <= 16'h0512;    16'd59891: out <= 16'hFF6B;
    16'd59892: out <= 16'h009F;    16'd59893: out <= 16'hF9A7;    16'd59894: out <= 16'h0666;    16'd59895: out <= 16'hFDB6;
    16'd59896: out <= 16'h0126;    16'd59897: out <= 16'hFACB;    16'd59898: out <= 16'h041E;    16'd59899: out <= 16'h06DA;
    16'd59900: out <= 16'hFF8F;    16'd59901: out <= 16'h018C;    16'd59902: out <= 16'h0289;    16'd59903: out <= 16'hF9B4;
    16'd59904: out <= 16'h0688;    16'd59905: out <= 16'h02CA;    16'd59906: out <= 16'h014D;    16'd59907: out <= 16'hFEE0;
    16'd59908: out <= 16'hFDA1;    16'd59909: out <= 16'h0764;    16'd59910: out <= 16'hFBAA;    16'd59911: out <= 16'hFEA8;
    16'd59912: out <= 16'h0396;    16'd59913: out <= 16'h0614;    16'd59914: out <= 16'hF902;    16'd59915: out <= 16'hFFDB;
    16'd59916: out <= 16'hFAF5;    16'd59917: out <= 16'hFFA5;    16'd59918: out <= 16'hFD2F;    16'd59919: out <= 16'h02F8;
    16'd59920: out <= 16'h0893;    16'd59921: out <= 16'h086A;    16'd59922: out <= 16'h0301;    16'd59923: out <= 16'hFAAE;
    16'd59924: out <= 16'h0483;    16'd59925: out <= 16'h0468;    16'd59926: out <= 16'h0677;    16'd59927: out <= 16'h02AA;
    16'd59928: out <= 16'hFCE3;    16'd59929: out <= 16'h035F;    16'd59930: out <= 16'h08C8;    16'd59931: out <= 16'hFE5E;
    16'd59932: out <= 16'hFAA7;    16'd59933: out <= 16'h0380;    16'd59934: out <= 16'hFF1B;    16'd59935: out <= 16'hFECA;
    16'd59936: out <= 16'hF9AE;    16'd59937: out <= 16'hFD03;    16'd59938: out <= 16'hFA81;    16'd59939: out <= 16'h019C;
    16'd59940: out <= 16'hFFC8;    16'd59941: out <= 16'hF852;    16'd59942: out <= 16'hFF02;    16'd59943: out <= 16'hF9A0;
    16'd59944: out <= 16'hFA4C;    16'd59945: out <= 16'hFE02;    16'd59946: out <= 16'h0136;    16'd59947: out <= 16'h0279;
    16'd59948: out <= 16'hFF3A;    16'd59949: out <= 16'h051C;    16'd59950: out <= 16'h04C9;    16'd59951: out <= 16'h059B;
    16'd59952: out <= 16'h0941;    16'd59953: out <= 16'h089E;    16'd59954: out <= 16'h0BAB;    16'd59955: out <= 16'h05CB;
    16'd59956: out <= 16'h08C6;    16'd59957: out <= 16'h02A2;    16'd59958: out <= 16'h0982;    16'd59959: out <= 16'hFB1F;
    16'd59960: out <= 16'h05EF;    16'd59961: out <= 16'h0010;    16'd59962: out <= 16'h07A1;    16'd59963: out <= 16'h0298;
    16'd59964: out <= 16'h011A;    16'd59965: out <= 16'h039F;    16'd59966: out <= 16'h062C;    16'd59967: out <= 16'h02D9;
    16'd59968: out <= 16'h0E41;    16'd59969: out <= 16'h0752;    16'd59970: out <= 16'h0B27;    16'd59971: out <= 16'h043A;
    16'd59972: out <= 16'h0061;    16'd59973: out <= 16'h0691;    16'd59974: out <= 16'h076B;    16'd59975: out <= 16'hFFF2;
    16'd59976: out <= 16'h0052;    16'd59977: out <= 16'hFF5A;    16'd59978: out <= 16'h07AC;    16'd59979: out <= 16'h044E;
    16'd59980: out <= 16'h0160;    16'd59981: out <= 16'h07BA;    16'd59982: out <= 16'h026B;    16'd59983: out <= 16'h0493;
    16'd59984: out <= 16'h04ED;    16'd59985: out <= 16'h08C3;    16'd59986: out <= 16'h0220;    16'd59987: out <= 16'hFFC3;
    16'd59988: out <= 16'h00A8;    16'd59989: out <= 16'h07DF;    16'd59990: out <= 16'hFE89;    16'd59991: out <= 16'hFF57;
    16'd59992: out <= 16'h0DA4;    16'd59993: out <= 16'hFF3A;    16'd59994: out <= 16'hFC23;    16'd59995: out <= 16'hFF44;
    16'd59996: out <= 16'h0005;    16'd59997: out <= 16'hFFD7;    16'd59998: out <= 16'hFBA4;    16'd59999: out <= 16'hFE2F;
    16'd60000: out <= 16'hFD94;    16'd60001: out <= 16'h0325;    16'd60002: out <= 16'hFFA2;    16'd60003: out <= 16'h0211;
    16'd60004: out <= 16'h00BC;    16'd60005: out <= 16'hFB30;    16'd60006: out <= 16'h00FF;    16'd60007: out <= 16'hFC47;
    16'd60008: out <= 16'h02B4;    16'd60009: out <= 16'hFD60;    16'd60010: out <= 16'hFDE1;    16'd60011: out <= 16'hFB54;
    16'd60012: out <= 16'h06B7;    16'd60013: out <= 16'h0386;    16'd60014: out <= 16'h00A9;    16'd60015: out <= 16'hFEEB;
    16'd60016: out <= 16'hFE0A;    16'd60017: out <= 16'h05FE;    16'd60018: out <= 16'hFF56;    16'd60019: out <= 16'hFEE8;
    16'd60020: out <= 16'h038B;    16'd60021: out <= 16'h014E;    16'd60022: out <= 16'hFF24;    16'd60023: out <= 16'h0457;
    16'd60024: out <= 16'hFF0A;    16'd60025: out <= 16'h00AA;    16'd60026: out <= 16'h0372;    16'd60027: out <= 16'h004C;
    16'd60028: out <= 16'hFA8D;    16'd60029: out <= 16'h0010;    16'd60030: out <= 16'h053A;    16'd60031: out <= 16'h0592;
    16'd60032: out <= 16'hFFF5;    16'd60033: out <= 16'h02E7;    16'd60034: out <= 16'h02F7;    16'd60035: out <= 16'h078D;
    16'd60036: out <= 16'h03A5;    16'd60037: out <= 16'h00F9;    16'd60038: out <= 16'h096E;    16'd60039: out <= 16'h029A;
    16'd60040: out <= 16'h0C10;    16'd60041: out <= 16'h0126;    16'd60042: out <= 16'h0298;    16'd60043: out <= 16'h091F;
    16'd60044: out <= 16'h0347;    16'd60045: out <= 16'h05B4;    16'd60046: out <= 16'h0662;    16'd60047: out <= 16'h01DF;
    16'd60048: out <= 16'hFEB5;    16'd60049: out <= 16'h04AF;    16'd60050: out <= 16'h0AF3;    16'd60051: out <= 16'h025C;
    16'd60052: out <= 16'h0A3D;    16'd60053: out <= 16'h062F;    16'd60054: out <= 16'hFF81;    16'd60055: out <= 16'h0410;
    16'd60056: out <= 16'h03FC;    16'd60057: out <= 16'h01C2;    16'd60058: out <= 16'h09D2;    16'd60059: out <= 16'hFD4C;
    16'd60060: out <= 16'hFFFE;    16'd60061: out <= 16'h05AD;    16'd60062: out <= 16'h0567;    16'd60063: out <= 16'h0526;
    16'd60064: out <= 16'h0337;    16'd60065: out <= 16'h0528;    16'd60066: out <= 16'h0492;    16'd60067: out <= 16'h00B3;
    16'd60068: out <= 16'h055D;    16'd60069: out <= 16'h0150;    16'd60070: out <= 16'h0A6D;    16'd60071: out <= 16'h0315;
    16'd60072: out <= 16'hFE66;    16'd60073: out <= 16'hFD38;    16'd60074: out <= 16'hF915;    16'd60075: out <= 16'hFF6A;
    16'd60076: out <= 16'h016E;    16'd60077: out <= 16'h00CF;    16'd60078: out <= 16'h015C;    16'd60079: out <= 16'hFD0E;
    16'd60080: out <= 16'h005F;    16'd60081: out <= 16'hFDBB;    16'd60082: out <= 16'h049F;    16'd60083: out <= 16'h02A5;
    16'd60084: out <= 16'h057F;    16'd60085: out <= 16'hFFE5;    16'd60086: out <= 16'h04AF;    16'd60087: out <= 16'h064B;
    16'd60088: out <= 16'h0325;    16'd60089: out <= 16'h00F7;    16'd60090: out <= 16'h0040;    16'd60091: out <= 16'h07B2;
    16'd60092: out <= 16'h01BA;    16'd60093: out <= 16'h0795;    16'd60094: out <= 16'h078B;    16'd60095: out <= 16'hFA9C;
    16'd60096: out <= 16'hFCF1;    16'd60097: out <= 16'h0474;    16'd60098: out <= 16'h0450;    16'd60099: out <= 16'hFFA6;
    16'd60100: out <= 16'hFDFC;    16'd60101: out <= 16'hF94E;    16'd60102: out <= 16'hFE3C;    16'd60103: out <= 16'h048D;
    16'd60104: out <= 16'h0472;    16'd60105: out <= 16'hFE48;    16'd60106: out <= 16'h0597;    16'd60107: out <= 16'hFF3F;
    16'd60108: out <= 16'hFB8F;    16'd60109: out <= 16'h0232;    16'd60110: out <= 16'hFF70;    16'd60111: out <= 16'hFFC4;
    16'd60112: out <= 16'hFE44;    16'd60113: out <= 16'h04C4;    16'd60114: out <= 16'h020E;    16'd60115: out <= 16'hFD3F;
    16'd60116: out <= 16'h0209;    16'd60117: out <= 16'h025F;    16'd60118: out <= 16'h0205;    16'd60119: out <= 16'h00B5;
    16'd60120: out <= 16'h00F2;    16'd60121: out <= 16'h0379;    16'd60122: out <= 16'hFDBC;    16'd60123: out <= 16'hFB07;
    16'd60124: out <= 16'h0350;    16'd60125: out <= 16'h06FA;    16'd60126: out <= 16'hFD89;    16'd60127: out <= 16'hFFD4;
    16'd60128: out <= 16'hFD3A;    16'd60129: out <= 16'h042D;    16'd60130: out <= 16'h0632;    16'd60131: out <= 16'hFFC5;
    16'd60132: out <= 16'hFF4F;    16'd60133: out <= 16'hFE13;    16'd60134: out <= 16'h02C2;    16'd60135: out <= 16'hF9F5;
    16'd60136: out <= 16'hFFC7;    16'd60137: out <= 16'hFF17;    16'd60138: out <= 16'h0286;    16'd60139: out <= 16'h036C;
    16'd60140: out <= 16'h0080;    16'd60141: out <= 16'h01EE;    16'd60142: out <= 16'h0149;    16'd60143: out <= 16'h02C9;
    16'd60144: out <= 16'h0326;    16'd60145: out <= 16'h05A8;    16'd60146: out <= 16'h0118;    16'd60147: out <= 16'h05EC;
    16'd60148: out <= 16'h03DD;    16'd60149: out <= 16'h032E;    16'd60150: out <= 16'h02F7;    16'd60151: out <= 16'h03DE;
    16'd60152: out <= 16'h0110;    16'd60153: out <= 16'hFA27;    16'd60154: out <= 16'hFB60;    16'd60155: out <= 16'hFF5E;
    16'd60156: out <= 16'h0125;    16'd60157: out <= 16'h0495;    16'd60158: out <= 16'hFDBE;    16'd60159: out <= 16'hFEE4;
    16'd60160: out <= 16'h0419;    16'd60161: out <= 16'h0265;    16'd60162: out <= 16'h0016;    16'd60163: out <= 16'hFFC1;
    16'd60164: out <= 16'hFD92;    16'd60165: out <= 16'h0189;    16'd60166: out <= 16'h0174;    16'd60167: out <= 16'h00D7;
    16'd60168: out <= 16'hFBC2;    16'd60169: out <= 16'hFBE6;    16'd60170: out <= 16'h05E4;    16'd60171: out <= 16'hF914;
    16'd60172: out <= 16'hFBAF;    16'd60173: out <= 16'h02B4;    16'd60174: out <= 16'hFC3C;    16'd60175: out <= 16'h0333;
    16'd60176: out <= 16'h006F;    16'd60177: out <= 16'hFAFD;    16'd60178: out <= 16'hFE2E;    16'd60179: out <= 16'hFE0B;
    16'd60180: out <= 16'h0137;    16'd60181: out <= 16'h04FF;    16'd60182: out <= 16'h0020;    16'd60183: out <= 16'h0486;
    16'd60184: out <= 16'hFFC6;    16'd60185: out <= 16'hFA97;    16'd60186: out <= 16'h01AC;    16'd60187: out <= 16'hFC71;
    16'd60188: out <= 16'hFC02;    16'd60189: out <= 16'h0596;    16'd60190: out <= 16'h022C;    16'd60191: out <= 16'hFD08;
    16'd60192: out <= 16'h0389;    16'd60193: out <= 16'h00AD;    16'd60194: out <= 16'hFD1A;    16'd60195: out <= 16'h01E9;
    16'd60196: out <= 16'hFD23;    16'd60197: out <= 16'h089E;    16'd60198: out <= 16'hFAB2;    16'd60199: out <= 16'h0363;
    16'd60200: out <= 16'h0619;    16'd60201: out <= 16'h0618;    16'd60202: out <= 16'h083C;    16'd60203: out <= 16'h0879;
    16'd60204: out <= 16'h08C8;    16'd60205: out <= 16'hF791;    16'd60206: out <= 16'h0664;    16'd60207: out <= 16'h05FE;
    16'd60208: out <= 16'h0337;    16'd60209: out <= 16'h0182;    16'd60210: out <= 16'hFB56;    16'd60211: out <= 16'h073F;
    16'd60212: out <= 16'h0C24;    16'd60213: out <= 16'h0210;    16'd60214: out <= 16'hFEDD;    16'd60215: out <= 16'h0A61;
    16'd60216: out <= 16'h06A8;    16'd60217: out <= 16'hFF3C;    16'd60218: out <= 16'h0529;    16'd60219: out <= 16'h0AD9;
    16'd60220: out <= 16'hFFC0;    16'd60221: out <= 16'hFBC4;    16'd60222: out <= 16'hF89A;    16'd60223: out <= 16'h037A;
    16'd60224: out <= 16'hFFA3;    16'd60225: out <= 16'h0614;    16'd60226: out <= 16'h02C0;    16'd60227: out <= 16'h045A;
    16'd60228: out <= 16'hFF67;    16'd60229: out <= 16'h01F0;    16'd60230: out <= 16'h0857;    16'd60231: out <= 16'hFD5B;
    16'd60232: out <= 16'h09B8;    16'd60233: out <= 16'hFFCE;    16'd60234: out <= 16'h004F;    16'd60235: out <= 16'h053C;
    16'd60236: out <= 16'h062A;    16'd60237: out <= 16'h05F6;    16'd60238: out <= 16'hFFBB;    16'd60239: out <= 16'h0091;
    16'd60240: out <= 16'hFF5F;    16'd60241: out <= 16'h0843;    16'd60242: out <= 16'h018B;    16'd60243: out <= 16'hFF67;
    16'd60244: out <= 16'h0A4F;    16'd60245: out <= 16'h0301;    16'd60246: out <= 16'h05AE;    16'd60247: out <= 16'h0AA9;
    16'd60248: out <= 16'h0B73;    16'd60249: out <= 16'h0314;    16'd60250: out <= 16'hFFA4;    16'd60251: out <= 16'hFD28;
    16'd60252: out <= 16'h03F3;    16'd60253: out <= 16'hFE55;    16'd60254: out <= 16'h06DC;    16'd60255: out <= 16'hFF5C;
    16'd60256: out <= 16'hFDA6;    16'd60257: out <= 16'h0127;    16'd60258: out <= 16'h00EA;    16'd60259: out <= 16'hFAE2;
    16'd60260: out <= 16'h0667;    16'd60261: out <= 16'hFE60;    16'd60262: out <= 16'hFEA9;    16'd60263: out <= 16'h03A7;
    16'd60264: out <= 16'hFE74;    16'd60265: out <= 16'h0715;    16'd60266: out <= 16'h0213;    16'd60267: out <= 16'hFAB0;
    16'd60268: out <= 16'hFB7D;    16'd60269: out <= 16'h02BD;    16'd60270: out <= 16'hFB1E;    16'd60271: out <= 16'hFF4C;
    16'd60272: out <= 16'hFC31;    16'd60273: out <= 16'h0075;    16'd60274: out <= 16'h0273;    16'd60275: out <= 16'h011F;
    16'd60276: out <= 16'hFDAB;    16'd60277: out <= 16'hFB5E;    16'd60278: out <= 16'hFD0F;    16'd60279: out <= 16'h036C;
    16'd60280: out <= 16'h0603;    16'd60281: out <= 16'h020D;    16'd60282: out <= 16'hFDF5;    16'd60283: out <= 16'hF2A6;
    16'd60284: out <= 16'hFEE5;    16'd60285: out <= 16'hFF79;    16'd60286: out <= 16'h0315;    16'd60287: out <= 16'hFC17;
    16'd60288: out <= 16'h01CB;    16'd60289: out <= 16'h0393;    16'd60290: out <= 16'h02E6;    16'd60291: out <= 16'h06FE;
    16'd60292: out <= 16'h020A;    16'd60293: out <= 16'h02D5;    16'd60294: out <= 16'h0333;    16'd60295: out <= 16'hFDD0;
    16'd60296: out <= 16'hFD8E;    16'd60297: out <= 16'h0579;    16'd60298: out <= 16'h0712;    16'd60299: out <= 16'h068A;
    16'd60300: out <= 16'hFF78;    16'd60301: out <= 16'h005A;    16'd60302: out <= 16'h03A6;    16'd60303: out <= 16'h0E19;
    16'd60304: out <= 16'h035E;    16'd60305: out <= 16'hFE80;    16'd60306: out <= 16'h0718;    16'd60307: out <= 16'h0227;
    16'd60308: out <= 16'h0A2A;    16'd60309: out <= 16'h0745;    16'd60310: out <= 16'h016E;    16'd60311: out <= 16'h076C;
    16'd60312: out <= 16'h052A;    16'd60313: out <= 16'h044D;    16'd60314: out <= 16'h0CB7;    16'd60315: out <= 16'h0B99;
    16'd60316: out <= 16'h0A18;    16'd60317: out <= 16'hF9DA;    16'd60318: out <= 16'h03B6;    16'd60319: out <= 16'h069B;
    16'd60320: out <= 16'h06F5;    16'd60321: out <= 16'hFF6E;    16'd60322: out <= 16'h0480;    16'd60323: out <= 16'hFB35;
    16'd60324: out <= 16'h02A7;    16'd60325: out <= 16'h0483;    16'd60326: out <= 16'hFE34;    16'd60327: out <= 16'hFBA4;
    16'd60328: out <= 16'hFE27;    16'd60329: out <= 16'h0297;    16'd60330: out <= 16'hF93F;    16'd60331: out <= 16'hFC59;
    16'd60332: out <= 16'h0510;    16'd60333: out <= 16'hFF7F;    16'd60334: out <= 16'h03BF;    16'd60335: out <= 16'h0750;
    16'd60336: out <= 16'hFE3C;    16'd60337: out <= 16'h0876;    16'd60338: out <= 16'h037A;    16'd60339: out <= 16'hFE9E;
    16'd60340: out <= 16'h0475;    16'd60341: out <= 16'hFB4F;    16'd60342: out <= 16'h0930;    16'd60343: out <= 16'h0590;
    16'd60344: out <= 16'h05A4;    16'd60345: out <= 16'h0A61;    16'd60346: out <= 16'h002E;    16'd60347: out <= 16'h0465;
    16'd60348: out <= 16'h0339;    16'd60349: out <= 16'hF983;    16'd60350: out <= 16'h05C1;    16'd60351: out <= 16'h03D5;
    16'd60352: out <= 16'h00A3;    16'd60353: out <= 16'hFFD8;    16'd60354: out <= 16'hFF61;    16'd60355: out <= 16'h06DD;
    16'd60356: out <= 16'hFBAA;    16'd60357: out <= 16'hFB51;    16'd60358: out <= 16'h00D2;    16'd60359: out <= 16'hFFAE;
    16'd60360: out <= 16'hF920;    16'd60361: out <= 16'h007F;    16'd60362: out <= 16'hFF16;    16'd60363: out <= 16'h029E;
    16'd60364: out <= 16'h0154;    16'd60365: out <= 16'hFEE0;    16'd60366: out <= 16'h076C;    16'd60367: out <= 16'h043C;
    16'd60368: out <= 16'h07A5;    16'd60369: out <= 16'h0205;    16'd60370: out <= 16'hFF62;    16'd60371: out <= 16'hF837;
    16'd60372: out <= 16'h0A5D;    16'd60373: out <= 16'h0268;    16'd60374: out <= 16'h017D;    16'd60375: out <= 16'hFC9E;
    16'd60376: out <= 16'hFE89;    16'd60377: out <= 16'hFCAF;    16'd60378: out <= 16'hFB3D;    16'd60379: out <= 16'hF8C6;
    16'd60380: out <= 16'h01A3;    16'd60381: out <= 16'hFDBB;    16'd60382: out <= 16'h0114;    16'd60383: out <= 16'h034C;
    16'd60384: out <= 16'h0026;    16'd60385: out <= 16'h088A;    16'd60386: out <= 16'h0301;    16'd60387: out <= 16'h0609;
    16'd60388: out <= 16'h03A4;    16'd60389: out <= 16'hFF1D;    16'd60390: out <= 16'h010B;    16'd60391: out <= 16'hFE20;
    16'd60392: out <= 16'h0AFB;    16'd60393: out <= 16'h01D8;    16'd60394: out <= 16'h0415;    16'd60395: out <= 16'hFE36;
    16'd60396: out <= 16'h02CC;    16'd60397: out <= 16'h0403;    16'd60398: out <= 16'h0340;    16'd60399: out <= 16'h0230;
    16'd60400: out <= 16'hFFAC;    16'd60401: out <= 16'h0070;    16'd60402: out <= 16'hFDE8;    16'd60403: out <= 16'h056F;
    16'd60404: out <= 16'h003D;    16'd60405: out <= 16'hFE14;    16'd60406: out <= 16'hFB94;    16'd60407: out <= 16'hFC4A;
    16'd60408: out <= 16'h046A;    16'd60409: out <= 16'h04F7;    16'd60410: out <= 16'h0074;    16'd60411: out <= 16'hFD0E;
    16'd60412: out <= 16'hF7A2;    16'd60413: out <= 16'hFB45;    16'd60414: out <= 16'h024D;    16'd60415: out <= 16'h0538;
    16'd60416: out <= 16'hFF9E;    16'd60417: out <= 16'h01A8;    16'd60418: out <= 16'h0363;    16'd60419: out <= 16'h03B1;
    16'd60420: out <= 16'h01BD;    16'd60421: out <= 16'hFFCD;    16'd60422: out <= 16'hFF66;    16'd60423: out <= 16'h011A;
    16'd60424: out <= 16'hFD53;    16'd60425: out <= 16'hFB8A;    16'd60426: out <= 16'h018D;    16'd60427: out <= 16'hFE5F;
    16'd60428: out <= 16'hFED2;    16'd60429: out <= 16'hFA7C;    16'd60430: out <= 16'h046F;    16'd60431: out <= 16'hFFD8;
    16'd60432: out <= 16'h0105;    16'd60433: out <= 16'hFE5C;    16'd60434: out <= 16'h0025;    16'd60435: out <= 16'hFF2C;
    16'd60436: out <= 16'hFD0B;    16'd60437: out <= 16'hFFCA;    16'd60438: out <= 16'h0257;    16'd60439: out <= 16'h01C7;
    16'd60440: out <= 16'h0054;    16'd60441: out <= 16'h026D;    16'd60442: out <= 16'hFBF4;    16'd60443: out <= 16'hFE22;
    16'd60444: out <= 16'h01D5;    16'd60445: out <= 16'h04CD;    16'd60446: out <= 16'hFF8D;    16'd60447: out <= 16'hFC0F;
    16'd60448: out <= 16'hFE5C;    16'd60449: out <= 16'hFF86;    16'd60450: out <= 16'hFCB1;    16'd60451: out <= 16'h06F6;
    16'd60452: out <= 16'h01B6;    16'd60453: out <= 16'h0558;    16'd60454: out <= 16'h03D4;    16'd60455: out <= 16'hFBB7;
    16'd60456: out <= 16'h002B;    16'd60457: out <= 16'hFF5F;    16'd60458: out <= 16'hFF8D;    16'd60459: out <= 16'hFD36;
    16'd60460: out <= 16'hFC32;    16'd60461: out <= 16'hF8C1;    16'd60462: out <= 16'h05DD;    16'd60463: out <= 16'h04C3;
    16'd60464: out <= 16'hFE6D;    16'd60465: out <= 16'h0A72;    16'd60466: out <= 16'h07AA;    16'd60467: out <= 16'h060D;
    16'd60468: out <= 16'h0417;    16'd60469: out <= 16'h0A00;    16'd60470: out <= 16'h09CF;    16'd60471: out <= 16'h0383;
    16'd60472: out <= 16'h0484;    16'd60473: out <= 16'h0509;    16'd60474: out <= 16'h0170;    16'd60475: out <= 16'h0916;
    16'd60476: out <= 16'h010A;    16'd60477: out <= 16'h06BD;    16'd60478: out <= 16'h062E;    16'd60479: out <= 16'h06FF;
    16'd60480: out <= 16'h036C;    16'd60481: out <= 16'h05D6;    16'd60482: out <= 16'h0022;    16'd60483: out <= 16'h090B;
    16'd60484: out <= 16'h031A;    16'd60485: out <= 16'h05AC;    16'd60486: out <= 16'h0DD4;    16'd60487: out <= 16'h0580;
    16'd60488: out <= 16'h03DA;    16'd60489: out <= 16'hFCD3;    16'd60490: out <= 16'h0195;    16'd60491: out <= 16'hFC8D;
    16'd60492: out <= 16'h075F;    16'd60493: out <= 16'hFCA3;    16'd60494: out <= 16'hFEA2;    16'd60495: out <= 16'h00B0;
    16'd60496: out <= 16'h0191;    16'd60497: out <= 16'h00B2;    16'd60498: out <= 16'h055B;    16'd60499: out <= 16'h0469;
    16'd60500: out <= 16'h02EC;    16'd60501: out <= 16'h00DB;    16'd60502: out <= 16'h0134;    16'd60503: out <= 16'h0810;
    16'd60504: out <= 16'hFA7D;    16'd60505: out <= 16'hFF08;    16'd60506: out <= 16'h009E;    16'd60507: out <= 16'hFEA2;
    16'd60508: out <= 16'hFD86;    16'd60509: out <= 16'hFFFC;    16'd60510: out <= 16'h003D;    16'd60511: out <= 16'hF957;
    16'd60512: out <= 16'hFD0E;    16'd60513: out <= 16'hFD9F;    16'd60514: out <= 16'hF46A;    16'd60515: out <= 16'h01BF;
    16'd60516: out <= 16'hFEB9;    16'd60517: out <= 16'h0425;    16'd60518: out <= 16'h0598;    16'd60519: out <= 16'h05CC;
    16'd60520: out <= 16'h01EA;    16'd60521: out <= 16'hFFE6;    16'd60522: out <= 16'h0261;    16'd60523: out <= 16'hFD63;
    16'd60524: out <= 16'h01AC;    16'd60525: out <= 16'hFFD4;    16'd60526: out <= 16'hFB57;    16'd60527: out <= 16'hFDAF;
    16'd60528: out <= 16'hFE47;    16'd60529: out <= 16'hFD9F;    16'd60530: out <= 16'h019E;    16'd60531: out <= 16'h041E;
    16'd60532: out <= 16'h043A;    16'd60533: out <= 16'hFF71;    16'd60534: out <= 16'hFCEF;    16'd60535: out <= 16'hFDC7;
    16'd60536: out <= 16'h04DE;    16'd60537: out <= 16'hFE5B;    16'd60538: out <= 16'h0A50;    16'd60539: out <= 16'h0411;
    16'd60540: out <= 16'h0344;    16'd60541: out <= 16'h0114;    16'd60542: out <= 16'hFC4B;    16'd60543: out <= 16'h0040;
    16'd60544: out <= 16'hFEC5;    16'd60545: out <= 16'hFB3C;    16'd60546: out <= 16'h0323;    16'd60547: out <= 16'h08DF;
    16'd60548: out <= 16'h01FE;    16'd60549: out <= 16'hFC27;    16'd60550: out <= 16'h00D9;    16'd60551: out <= 16'h09E0;
    16'd60552: out <= 16'h0534;    16'd60553: out <= 16'h06F6;    16'd60554: out <= 16'h0469;    16'd60555: out <= 16'hFA31;
    16'd60556: out <= 16'hFDD2;    16'd60557: out <= 16'h0607;    16'd60558: out <= 16'h00BA;    16'd60559: out <= 16'h07EC;
    16'd60560: out <= 16'hFE55;    16'd60561: out <= 16'h068E;    16'd60562: out <= 16'h01CF;    16'd60563: out <= 16'h003E;
    16'd60564: out <= 16'h002B;    16'd60565: out <= 16'h03E9;    16'd60566: out <= 16'h06A2;    16'd60567: out <= 16'h0270;
    16'd60568: out <= 16'h0614;    16'd60569: out <= 16'h0078;    16'd60570: out <= 16'h0993;    16'd60571: out <= 16'h0314;
    16'd60572: out <= 16'h0181;    16'd60573: out <= 16'h053C;    16'd60574: out <= 16'hF8BE;    16'd60575: out <= 16'h03CF;
    16'd60576: out <= 16'h004A;    16'd60577: out <= 16'hFFD5;    16'd60578: out <= 16'h0B15;    16'd60579: out <= 16'h0388;
    16'd60580: out <= 16'h0300;    16'd60581: out <= 16'hFAB5;    16'd60582: out <= 16'hFC04;    16'd60583: out <= 16'h0133;
    16'd60584: out <= 16'hFF9D;    16'd60585: out <= 16'hFFE5;    16'd60586: out <= 16'h017A;    16'd60587: out <= 16'hF9E2;
    16'd60588: out <= 16'h03F2;    16'd60589: out <= 16'hFEDD;    16'd60590: out <= 16'hF2DB;    16'd60591: out <= 16'h097E;
    16'd60592: out <= 16'hFFFB;    16'd60593: out <= 16'h03F5;    16'd60594: out <= 16'h0394;    16'd60595: out <= 16'h0D5B;
    16'd60596: out <= 16'h03B5;    16'd60597: out <= 16'hFB52;    16'd60598: out <= 16'h02EB;    16'd60599: out <= 16'hFD5A;
    16'd60600: out <= 16'hFE5E;    16'd60601: out <= 16'h005C;    16'd60602: out <= 16'h0136;    16'd60603: out <= 16'hFEF6;
    16'd60604: out <= 16'h01AB;    16'd60605: out <= 16'h0142;    16'd60606: out <= 16'h01FC;    16'd60607: out <= 16'h0312;
    16'd60608: out <= 16'hF87E;    16'd60609: out <= 16'h01A8;    16'd60610: out <= 16'h0441;    16'd60611: out <= 16'h028C;
    16'd60612: out <= 16'hFAB3;    16'd60613: out <= 16'hF9C4;    16'd60614: out <= 16'hFBD3;    16'd60615: out <= 16'hFEBB;
    16'd60616: out <= 16'hFB90;    16'd60617: out <= 16'h004A;    16'd60618: out <= 16'hF9A1;    16'd60619: out <= 16'hF52E;
    16'd60620: out <= 16'h023E;    16'd60621: out <= 16'h05B3;    16'd60622: out <= 16'h0115;    16'd60623: out <= 16'hFF77;
    16'd60624: out <= 16'h031E;    16'd60625: out <= 16'hFCE7;    16'd60626: out <= 16'hF90C;    16'd60627: out <= 16'h05AF;
    16'd60628: out <= 16'h0036;    16'd60629: out <= 16'hFAD9;    16'd60630: out <= 16'h0659;    16'd60631: out <= 16'hFEE3;
    16'd60632: out <= 16'h00F3;    16'd60633: out <= 16'h01DB;    16'd60634: out <= 16'hFD5C;    16'd60635: out <= 16'hFEA6;
    16'd60636: out <= 16'h03BB;    16'd60637: out <= 16'hFF8E;    16'd60638: out <= 16'hFFEA;    16'd60639: out <= 16'hFA42;
    16'd60640: out <= 16'hF9D5;    16'd60641: out <= 16'h0151;    16'd60642: out <= 16'h017A;    16'd60643: out <= 16'hFF72;
    16'd60644: out <= 16'h07FF;    16'd60645: out <= 16'h0097;    16'd60646: out <= 16'h009E;    16'd60647: out <= 16'h031C;
    16'd60648: out <= 16'hFEA4;    16'd60649: out <= 16'h070F;    16'd60650: out <= 16'h017F;    16'd60651: out <= 16'h082E;
    16'd60652: out <= 16'hF766;    16'd60653: out <= 16'hFA9C;    16'd60654: out <= 16'h0270;    16'd60655: out <= 16'hFD9B;
    16'd60656: out <= 16'h0152;    16'd60657: out <= 16'h002F;    16'd60658: out <= 16'hFFD6;    16'd60659: out <= 16'h05B3;
    16'd60660: out <= 16'hF989;    16'd60661: out <= 16'hFE26;    16'd60662: out <= 16'hFB8C;    16'd60663: out <= 16'hFD83;
    16'd60664: out <= 16'hFA4C;    16'd60665: out <= 16'hFCD3;    16'd60666: out <= 16'h00A3;    16'd60667: out <= 16'hFED4;
    16'd60668: out <= 16'hFCFB;    16'd60669: out <= 16'hFEF6;    16'd60670: out <= 16'h0204;    16'd60671: out <= 16'hFC22;
    16'd60672: out <= 16'hF9CD;    16'd60673: out <= 16'hFF9D;    16'd60674: out <= 16'hFF15;    16'd60675: out <= 16'hF91D;
    16'd60676: out <= 16'hFF12;    16'd60677: out <= 16'h0040;    16'd60678: out <= 16'hFE5D;    16'd60679: out <= 16'hFC06;
    16'd60680: out <= 16'h0195;    16'd60681: out <= 16'h02BC;    16'd60682: out <= 16'h05EA;    16'd60683: out <= 16'h0169;
    16'd60684: out <= 16'h01C2;    16'd60685: out <= 16'h0735;    16'd60686: out <= 16'h04C0;    16'd60687: out <= 16'hFD82;
    16'd60688: out <= 16'hFFC9;    16'd60689: out <= 16'h01A7;    16'd60690: out <= 16'hFE47;    16'd60691: out <= 16'hFD10;
    16'd60692: out <= 16'hF60A;    16'd60693: out <= 16'hFF16;    16'd60694: out <= 16'h0200;    16'd60695: out <= 16'hFE31;
    16'd60696: out <= 16'h0492;    16'd60697: out <= 16'hF8C4;    16'd60698: out <= 16'hFD49;    16'd60699: out <= 16'h000F;
    16'd60700: out <= 16'hFD9C;    16'd60701: out <= 16'hFBB3;    16'd60702: out <= 16'h0570;    16'd60703: out <= 16'h03E4;
    16'd60704: out <= 16'hFFBA;    16'd60705: out <= 16'h02F6;    16'd60706: out <= 16'hFC0C;    16'd60707: out <= 16'hFCF1;
    16'd60708: out <= 16'hFC5F;    16'd60709: out <= 16'hFFA4;    16'd60710: out <= 16'hFF17;    16'd60711: out <= 16'h01C7;
    16'd60712: out <= 16'hFE15;    16'd60713: out <= 16'h006B;    16'd60714: out <= 16'hFF55;    16'd60715: out <= 16'h06B4;
    16'd60716: out <= 16'h03EC;    16'd60717: out <= 16'hFFF1;    16'd60718: out <= 16'h068F;    16'd60719: out <= 16'h0225;
    16'd60720: out <= 16'h0460;    16'd60721: out <= 16'h09D1;    16'd60722: out <= 16'h071E;    16'd60723: out <= 16'h056F;
    16'd60724: out <= 16'h0143;    16'd60725: out <= 16'h0721;    16'd60726: out <= 16'h05FD;    16'd60727: out <= 16'h005F;
    16'd60728: out <= 16'h016C;    16'd60729: out <= 16'h04EA;    16'd60730: out <= 16'h03EE;    16'd60731: out <= 16'h0122;
    16'd60732: out <= 16'h021D;    16'd60733: out <= 16'h035E;    16'd60734: out <= 16'h04D8;    16'd60735: out <= 16'h01A2;
    16'd60736: out <= 16'h0057;    16'd60737: out <= 16'h01F8;    16'd60738: out <= 16'h057E;    16'd60739: out <= 16'hFDA5;
    16'd60740: out <= 16'h0BEC;    16'd60741: out <= 16'h0163;    16'd60742: out <= 16'hFFE0;    16'd60743: out <= 16'h0289;
    16'd60744: out <= 16'h00A9;    16'd60745: out <= 16'h07F5;    16'd60746: out <= 16'h0365;    16'd60747: out <= 16'h03A7;
    16'd60748: out <= 16'h03E7;    16'd60749: out <= 16'h0043;    16'd60750: out <= 16'h0252;    16'd60751: out <= 16'h078A;
    16'd60752: out <= 16'h01F2;    16'd60753: out <= 16'h01BA;    16'd60754: out <= 16'h02FE;    16'd60755: out <= 16'h0566;
    16'd60756: out <= 16'h0448;    16'd60757: out <= 16'h06D9;    16'd60758: out <= 16'h013A;    16'd60759: out <= 16'hFFD5;
    16'd60760: out <= 16'h025C;    16'd60761: out <= 16'hFD35;    16'd60762: out <= 16'hFB73;    16'd60763: out <= 16'h04AA;
    16'd60764: out <= 16'h00E5;    16'd60765: out <= 16'h0241;    16'd60766: out <= 16'h00E6;    16'd60767: out <= 16'h039A;
    16'd60768: out <= 16'h01D9;    16'd60769: out <= 16'h0253;    16'd60770: out <= 16'hFB55;    16'd60771: out <= 16'hFF5B;
    16'd60772: out <= 16'h084C;    16'd60773: out <= 16'h0358;    16'd60774: out <= 16'hFB9D;    16'd60775: out <= 16'h0107;
    16'd60776: out <= 16'h01A6;    16'd60777: out <= 16'hFCCB;    16'd60778: out <= 16'hFD00;    16'd60779: out <= 16'h0982;
    16'd60780: out <= 16'hFB75;    16'd60781: out <= 16'h0295;    16'd60782: out <= 16'hFD98;    16'd60783: out <= 16'h062B;
    16'd60784: out <= 16'hFAF0;    16'd60785: out <= 16'hFF8E;    16'd60786: out <= 16'h0235;    16'd60787: out <= 16'hFA11;
    16'd60788: out <= 16'hFBC7;    16'd60789: out <= 16'hFFCA;    16'd60790: out <= 16'hFADA;    16'd60791: out <= 16'h025F;
    16'd60792: out <= 16'hFF89;    16'd60793: out <= 16'h0A94;    16'd60794: out <= 16'h06A7;    16'd60795: out <= 16'h04A4;
    16'd60796: out <= 16'h0556;    16'd60797: out <= 16'hF785;    16'd60798: out <= 16'h03AE;    16'd60799: out <= 16'hFEBC;
    16'd60800: out <= 16'hFB2E;    16'd60801: out <= 16'h00D3;    16'd60802: out <= 16'hF8D5;    16'd60803: out <= 16'h026C;
    16'd60804: out <= 16'hFDAB;    16'd60805: out <= 16'h0295;    16'd60806: out <= 16'h050E;    16'd60807: out <= 16'hFE4A;
    16'd60808: out <= 16'h044A;    16'd60809: out <= 16'h024D;    16'd60810: out <= 16'hFD2B;    16'd60811: out <= 16'h0009;
    16'd60812: out <= 16'h046B;    16'd60813: out <= 16'h065E;    16'd60814: out <= 16'h038B;    16'd60815: out <= 16'h05B7;
    16'd60816: out <= 16'h0AC7;    16'd60817: out <= 16'hFF34;    16'd60818: out <= 16'h0017;    16'd60819: out <= 16'h0112;
    16'd60820: out <= 16'h037E;    16'd60821: out <= 16'h00F3;    16'd60822: out <= 16'h041B;    16'd60823: out <= 16'h071D;
    16'd60824: out <= 16'hFF43;    16'd60825: out <= 16'hFD7A;    16'd60826: out <= 16'h0335;    16'd60827: out <= 16'h044F;
    16'd60828: out <= 16'hFB8E;    16'd60829: out <= 16'hFA3F;    16'd60830: out <= 16'hFF65;    16'd60831: out <= 16'h07BA;
    16'd60832: out <= 16'hFFEE;    16'd60833: out <= 16'h05BC;    16'd60834: out <= 16'h00B0;    16'd60835: out <= 16'h02A2;
    16'd60836: out <= 16'h048D;    16'd60837: out <= 16'h01F3;    16'd60838: out <= 16'hFCB9;    16'd60839: out <= 16'hFE16;
    16'd60840: out <= 16'h00EE;    16'd60841: out <= 16'h0473;    16'd60842: out <= 16'hFE5B;    16'd60843: out <= 16'h0556;
    16'd60844: out <= 16'h031C;    16'd60845: out <= 16'h023F;    16'd60846: out <= 16'h0969;    16'd60847: out <= 16'h00DA;
    16'd60848: out <= 16'h0023;    16'd60849: out <= 16'h04E8;    16'd60850: out <= 16'h01CF;    16'd60851: out <= 16'h0806;
    16'd60852: out <= 16'h0780;    16'd60853: out <= 16'h0120;    16'd60854: out <= 16'h009B;    16'd60855: out <= 16'h01CC;
    16'd60856: out <= 16'h0006;    16'd60857: out <= 16'h097B;    16'd60858: out <= 16'h0806;    16'd60859: out <= 16'h06F7;
    16'd60860: out <= 16'hFCFD;    16'd60861: out <= 16'hFE5A;    16'd60862: out <= 16'h0388;    16'd60863: out <= 16'h0416;
    16'd60864: out <= 16'h045C;    16'd60865: out <= 16'hFD30;    16'd60866: out <= 16'h04A1;    16'd60867: out <= 16'h042C;
    16'd60868: out <= 16'h043D;    16'd60869: out <= 16'h0503;    16'd60870: out <= 16'hFE2E;    16'd60871: out <= 16'h0305;
    16'd60872: out <= 16'hF98A;    16'd60873: out <= 16'hF9F2;    16'd60874: out <= 16'h0093;    16'd60875: out <= 16'hF9AE;
    16'd60876: out <= 16'h0359;    16'd60877: out <= 16'hFC1B;    16'd60878: out <= 16'h0991;    16'd60879: out <= 16'h0338;
    16'd60880: out <= 16'hFB58;    16'd60881: out <= 16'h04FE;    16'd60882: out <= 16'h04DF;    16'd60883: out <= 16'hFF62;
    16'd60884: out <= 16'h03C1;    16'd60885: out <= 16'h0068;    16'd60886: out <= 16'h0756;    16'd60887: out <= 16'h0606;
    16'd60888: out <= 16'h050E;    16'd60889: out <= 16'hFE17;    16'd60890: out <= 16'hF829;    16'd60891: out <= 16'hFF18;
    16'd60892: out <= 16'hFFC8;    16'd60893: out <= 16'hFF9A;    16'd60894: out <= 16'h034B;    16'd60895: out <= 16'hFDF1;
    16'd60896: out <= 16'hFC66;    16'd60897: out <= 16'hFEE2;    16'd60898: out <= 16'h021E;    16'd60899: out <= 16'hFECD;
    16'd60900: out <= 16'h00EF;    16'd60901: out <= 16'hFB59;    16'd60902: out <= 16'hFE67;    16'd60903: out <= 16'h0146;
    16'd60904: out <= 16'h0073;    16'd60905: out <= 16'hFF38;    16'd60906: out <= 16'hFB0E;    16'd60907: out <= 16'h0101;
    16'd60908: out <= 16'hFD57;    16'd60909: out <= 16'h0563;    16'd60910: out <= 16'h023D;    16'd60911: out <= 16'h027A;
    16'd60912: out <= 16'hFE1B;    16'd60913: out <= 16'hFF97;    16'd60914: out <= 16'hFC20;    16'd60915: out <= 16'h0634;
    16'd60916: out <= 16'hFECE;    16'd60917: out <= 16'h00D4;    16'd60918: out <= 16'hFA43;    16'd60919: out <= 16'h048C;
    16'd60920: out <= 16'hFC81;    16'd60921: out <= 16'h00D6;    16'd60922: out <= 16'hFD74;    16'd60923: out <= 16'h0050;
    16'd60924: out <= 16'hFB02;    16'd60925: out <= 16'hFED7;    16'd60926: out <= 16'h06D5;    16'd60927: out <= 16'hFF34;
    16'd60928: out <= 16'h0536;    16'd60929: out <= 16'hFF70;    16'd60930: out <= 16'hFABB;    16'd60931: out <= 16'hF712;
    16'd60932: out <= 16'h01CD;    16'd60933: out <= 16'h0663;    16'd60934: out <= 16'hFA4F;    16'd60935: out <= 16'hFCFE;
    16'd60936: out <= 16'h04D7;    16'd60937: out <= 16'h03DF;    16'd60938: out <= 16'h0277;    16'd60939: out <= 16'hFF76;
    16'd60940: out <= 16'hFCDD;    16'd60941: out <= 16'h0125;    16'd60942: out <= 16'h0522;    16'd60943: out <= 16'hFBC5;
    16'd60944: out <= 16'h0100;    16'd60945: out <= 16'h0340;    16'd60946: out <= 16'hFD53;    16'd60947: out <= 16'hFC72;
    16'd60948: out <= 16'h0199;    16'd60949: out <= 16'h0891;    16'd60950: out <= 16'hFCE0;    16'd60951: out <= 16'hFE10;
    16'd60952: out <= 16'hF837;    16'd60953: out <= 16'h076F;    16'd60954: out <= 16'h0212;    16'd60955: out <= 16'hFF8A;
    16'd60956: out <= 16'hFBEC;    16'd60957: out <= 16'h026A;    16'd60958: out <= 16'h0486;    16'd60959: out <= 16'hFF27;
    16'd60960: out <= 16'hF941;    16'd60961: out <= 16'h0284;    16'd60962: out <= 16'h041A;    16'd60963: out <= 16'h01CC;
    16'd60964: out <= 16'hFED9;    16'd60965: out <= 16'hFD01;    16'd60966: out <= 16'h00B4;    16'd60967: out <= 16'hF80D;
    16'd60968: out <= 16'h0262;    16'd60969: out <= 16'h0335;    16'd60970: out <= 16'h017B;    16'd60971: out <= 16'hFD61;
    16'd60972: out <= 16'h04D9;    16'd60973: out <= 16'hFE6C;    16'd60974: out <= 16'h0440;    16'd60975: out <= 16'h01A3;
    16'd60976: out <= 16'h0CF0;    16'd60977: out <= 16'h02D1;    16'd60978: out <= 16'h0568;    16'd60979: out <= 16'h0143;
    16'd60980: out <= 16'h026E;    16'd60981: out <= 16'h0425;    16'd60982: out <= 16'h0387;    16'd60983: out <= 16'h07B1;
    16'd60984: out <= 16'h0424;    16'd60985: out <= 16'h053A;    16'd60986: out <= 16'h01F0;    16'd60987: out <= 16'h05C2;
    16'd60988: out <= 16'h005C;    16'd60989: out <= 16'h0488;    16'd60990: out <= 16'hFFD9;    16'd60991: out <= 16'h0354;
    16'd60992: out <= 16'h00E3;    16'd60993: out <= 16'hFFAE;    16'd60994: out <= 16'h04A1;    16'd60995: out <= 16'h06EC;
    16'd60996: out <= 16'h03EC;    16'd60997: out <= 16'h0086;    16'd60998: out <= 16'h0185;    16'd60999: out <= 16'h096F;
    16'd61000: out <= 16'h05AA;    16'd61001: out <= 16'h0241;    16'd61002: out <= 16'h005C;    16'd61003: out <= 16'h060E;
    16'd61004: out <= 16'hFC7E;    16'd61005: out <= 16'h03C1;    16'd61006: out <= 16'h0EFE;    16'd61007: out <= 16'h03AC;
    16'd61008: out <= 16'h01B8;    16'd61009: out <= 16'hFD03;    16'd61010: out <= 16'h0862;    16'd61011: out <= 16'hFF1C;
    16'd61012: out <= 16'hFC9C;    16'd61013: out <= 16'hFEE1;    16'd61014: out <= 16'h0300;    16'd61015: out <= 16'h065C;
    16'd61016: out <= 16'hFF6F;    16'd61017: out <= 16'hFD9F;    16'd61018: out <= 16'hFA19;    16'd61019: out <= 16'hFA6D;
    16'd61020: out <= 16'hFFEC;    16'd61021: out <= 16'h057B;    16'd61022: out <= 16'hFC99;    16'd61023: out <= 16'hFADF;
    16'd61024: out <= 16'h0207;    16'd61025: out <= 16'hFEE8;    16'd61026: out <= 16'h00A3;    16'd61027: out <= 16'h0B99;
    16'd61028: out <= 16'h06F7;    16'd61029: out <= 16'hFD02;    16'd61030: out <= 16'hFE18;    16'd61031: out <= 16'hFFEC;
    16'd61032: out <= 16'h0218;    16'd61033: out <= 16'hFF76;    16'd61034: out <= 16'hFFC3;    16'd61035: out <= 16'h009B;
    16'd61036: out <= 16'hFE34;    16'd61037: out <= 16'hFA45;    16'd61038: out <= 16'h0122;    16'd61039: out <= 16'h0314;
    16'd61040: out <= 16'h036C;    16'd61041: out <= 16'hFEF8;    16'd61042: out <= 16'h006F;    16'd61043: out <= 16'h0428;
    16'd61044: out <= 16'hFEB1;    16'd61045: out <= 16'h0537;    16'd61046: out <= 16'hFF30;    16'd61047: out <= 16'hFA5B;
    16'd61048: out <= 16'h01B8;    16'd61049: out <= 16'h045C;    16'd61050: out <= 16'hFF50;    16'd61051: out <= 16'hFA43;
    16'd61052: out <= 16'h018B;    16'd61053: out <= 16'hF9FC;    16'd61054: out <= 16'hFE6B;    16'd61055: out <= 16'hFCE4;
    16'd61056: out <= 16'hFF30;    16'd61057: out <= 16'h04C0;    16'd61058: out <= 16'h054F;    16'd61059: out <= 16'hFCA9;
    16'd61060: out <= 16'h0189;    16'd61061: out <= 16'h018E;    16'd61062: out <= 16'hFE89;    16'd61063: out <= 16'h041E;
    16'd61064: out <= 16'h024C;    16'd61065: out <= 16'h0174;    16'd61066: out <= 16'hFEC8;    16'd61067: out <= 16'h0181;
    16'd61068: out <= 16'hFD77;    16'd61069: out <= 16'hFAF4;    16'd61070: out <= 16'h0320;    16'd61071: out <= 16'hF514;
    16'd61072: out <= 16'h0144;    16'd61073: out <= 16'h0925;    16'd61074: out <= 16'h03C9;    16'd61075: out <= 16'hFE83;
    16'd61076: out <= 16'hFB60;    16'd61077: out <= 16'h0920;    16'd61078: out <= 16'h0162;    16'd61079: out <= 16'h0002;
    16'd61080: out <= 16'h00ED;    16'd61081: out <= 16'hFE9F;    16'd61082: out <= 16'h0180;    16'd61083: out <= 16'hFF5C;
    16'd61084: out <= 16'h02AB;    16'd61085: out <= 16'hFCDC;    16'd61086: out <= 16'h0112;    16'd61087: out <= 16'h02FF;
    16'd61088: out <= 16'hFCA8;    16'd61089: out <= 16'h015C;    16'd61090: out <= 16'h00AE;    16'd61091: out <= 16'h050A;
    16'd61092: out <= 16'hFA51;    16'd61093: out <= 16'hFC62;    16'd61094: out <= 16'h002A;    16'd61095: out <= 16'hFB13;
    16'd61096: out <= 16'hF8F7;    16'd61097: out <= 16'hFF46;    16'd61098: out <= 16'hFFE6;    16'd61099: out <= 16'hFF6B;
    16'd61100: out <= 16'h0543;    16'd61101: out <= 16'h0325;    16'd61102: out <= 16'h0918;    16'd61103: out <= 16'hFDD0;
    16'd61104: out <= 16'h0800;    16'd61105: out <= 16'h03D8;    16'd61106: out <= 16'h03F6;    16'd61107: out <= 16'h0211;
    16'd61108: out <= 16'h037C;    16'd61109: out <= 16'h034E;    16'd61110: out <= 16'h03E2;    16'd61111: out <= 16'h03CE;
    16'd61112: out <= 16'h0777;    16'd61113: out <= 16'h04B8;    16'd61114: out <= 16'h0009;    16'd61115: out <= 16'h0442;
    16'd61116: out <= 16'hFD4C;    16'd61117: out <= 16'h03A3;    16'd61118: out <= 16'h035F;    16'd61119: out <= 16'h038F;
    16'd61120: out <= 16'h035B;    16'd61121: out <= 16'h07ED;    16'd61122: out <= 16'h0492;    16'd61123: out <= 16'h00DC;
    16'd61124: out <= 16'hFED4;    16'd61125: out <= 16'hFE9E;    16'd61126: out <= 16'h0139;    16'd61127: out <= 16'h0612;
    16'd61128: out <= 16'h03F7;    16'd61129: out <= 16'h023C;    16'd61130: out <= 16'h0560;    16'd61131: out <= 16'h0137;
    16'd61132: out <= 16'hF852;    16'd61133: out <= 16'hFB2A;    16'd61134: out <= 16'h069C;    16'd61135: out <= 16'hFA0C;
    16'd61136: out <= 16'hFF9D;    16'd61137: out <= 16'hF80B;    16'd61138: out <= 16'hFE52;    16'd61139: out <= 16'hFCE6;
    16'd61140: out <= 16'hFDC7;    16'd61141: out <= 16'hFD77;    16'd61142: out <= 16'h0543;    16'd61143: out <= 16'h0133;
    16'd61144: out <= 16'hF78B;    16'd61145: out <= 16'hFDC8;    16'd61146: out <= 16'h00B3;    16'd61147: out <= 16'hFDC2;
    16'd61148: out <= 16'hFEAB;    16'd61149: out <= 16'hFF10;    16'd61150: out <= 16'hFAF0;    16'd61151: out <= 16'hFF9F;
    16'd61152: out <= 16'h0080;    16'd61153: out <= 16'hFE6A;    16'd61154: out <= 16'h009B;    16'd61155: out <= 16'h011B;
    16'd61156: out <= 16'hFDE8;    16'd61157: out <= 16'hFC69;    16'd61158: out <= 16'hFD0E;    16'd61159: out <= 16'h0017;
    16'd61160: out <= 16'h0282;    16'd61161: out <= 16'hFE67;    16'd61162: out <= 16'h01F9;    16'd61163: out <= 16'hF974;
    16'd61164: out <= 16'h0369;    16'd61165: out <= 16'hFF92;    16'd61166: out <= 16'hFD2B;    16'd61167: out <= 16'hF91E;
    16'd61168: out <= 16'hFC8B;    16'd61169: out <= 16'h02E5;    16'd61170: out <= 16'h013D;    16'd61171: out <= 16'hFECA;
    16'd61172: out <= 16'h0295;    16'd61173: out <= 16'h02C8;    16'd61174: out <= 16'hFDC3;    16'd61175: out <= 16'hFF29;
    16'd61176: out <= 16'h0453;    16'd61177: out <= 16'h051E;    16'd61178: out <= 16'hFB65;    16'd61179: out <= 16'h0382;
    16'd61180: out <= 16'h038C;    16'd61181: out <= 16'h0174;    16'd61182: out <= 16'h014A;    16'd61183: out <= 16'h0248;
    16'd61184: out <= 16'h0039;    16'd61185: out <= 16'h0569;    16'd61186: out <= 16'hF784;    16'd61187: out <= 16'h05F9;
    16'd61188: out <= 16'h0301;    16'd61189: out <= 16'hFFEA;    16'd61190: out <= 16'h046A;    16'd61191: out <= 16'h043E;
    16'd61192: out <= 16'h02E7;    16'd61193: out <= 16'h0053;    16'd61194: out <= 16'hFB02;    16'd61195: out <= 16'hFD76;
    16'd61196: out <= 16'hFE94;    16'd61197: out <= 16'hFEC4;    16'd61198: out <= 16'hFCE2;    16'd61199: out <= 16'hFB1F;
    16'd61200: out <= 16'hFFF7;    16'd61201: out <= 16'h02D6;    16'd61202: out <= 16'hFEA6;    16'd61203: out <= 16'hFB8B;
    16'd61204: out <= 16'h0175;    16'd61205: out <= 16'hFDD3;    16'd61206: out <= 16'h00BC;    16'd61207: out <= 16'h0168;
    16'd61208: out <= 16'hFECC;    16'd61209: out <= 16'h0382;    16'd61210: out <= 16'h06D0;    16'd61211: out <= 16'hFDB8;
    16'd61212: out <= 16'h04A4;    16'd61213: out <= 16'h020B;    16'd61214: out <= 16'h0026;    16'd61215: out <= 16'hFA93;
    16'd61216: out <= 16'h0291;    16'd61217: out <= 16'hFBB3;    16'd61218: out <= 16'hFE76;    16'd61219: out <= 16'h01DD;
    16'd61220: out <= 16'hFB6D;    16'd61221: out <= 16'hFFF8;    16'd61222: out <= 16'hFA55;    16'd61223: out <= 16'h0069;
    16'd61224: out <= 16'h02BF;    16'd61225: out <= 16'hFF56;    16'd61226: out <= 16'hF7C2;    16'd61227: out <= 16'h0134;
    16'd61228: out <= 16'h03F6;    16'd61229: out <= 16'h0568;    16'd61230: out <= 16'hFB9D;    16'd61231: out <= 16'h0781;
    16'd61232: out <= 16'h0739;    16'd61233: out <= 16'hFF47;    16'd61234: out <= 16'h0C78;    16'd61235: out <= 16'h04B9;
    16'd61236: out <= 16'hFBB7;    16'd61237: out <= 16'h0C72;    16'd61238: out <= 16'h0779;    16'd61239: out <= 16'h04C8;
    16'd61240: out <= 16'hFD1A;    16'd61241: out <= 16'h0552;    16'd61242: out <= 16'h030A;    16'd61243: out <= 16'h0241;
    16'd61244: out <= 16'h0AB4;    16'd61245: out <= 16'h04D1;    16'd61246: out <= 16'h0641;    16'd61247: out <= 16'h05E1;
    16'd61248: out <= 16'h0040;    16'd61249: out <= 16'h05B6;    16'd61250: out <= 16'h0771;    16'd61251: out <= 16'h0648;
    16'd61252: out <= 16'h0383;    16'd61253: out <= 16'h0142;    16'd61254: out <= 16'hFFB2;    16'd61255: out <= 16'hFD98;
    16'd61256: out <= 16'h0586;    16'd61257: out <= 16'h00D4;    16'd61258: out <= 16'h03EE;    16'd61259: out <= 16'h05EA;
    16'd61260: out <= 16'hFF7E;    16'd61261: out <= 16'h004C;    16'd61262: out <= 16'h02EF;    16'd61263: out <= 16'h08E0;
    16'd61264: out <= 16'h0464;    16'd61265: out <= 16'h06A3;    16'd61266: out <= 16'h0232;    16'd61267: out <= 16'hFEF0;
    16'd61268: out <= 16'hFD60;    16'd61269: out <= 16'hFF11;    16'd61270: out <= 16'hFF49;    16'd61271: out <= 16'hFF9C;
    16'd61272: out <= 16'h026C;    16'd61273: out <= 16'h0276;    16'd61274: out <= 16'hFC88;    16'd61275: out <= 16'hFC17;
    16'd61276: out <= 16'hF929;    16'd61277: out <= 16'h0302;    16'd61278: out <= 16'h047A;    16'd61279: out <= 16'h001D;
    16'd61280: out <= 16'hFCD8;    16'd61281: out <= 16'h07B1;    16'd61282: out <= 16'h01D7;    16'd61283: out <= 16'h02C0;
    16'd61284: out <= 16'hFEE6;    16'd61285: out <= 16'h00A9;    16'd61286: out <= 16'hFF50;    16'd61287: out <= 16'h0195;
    16'd61288: out <= 16'hFBAF;    16'd61289: out <= 16'h02D0;    16'd61290: out <= 16'h058D;    16'd61291: out <= 16'h003F;
    16'd61292: out <= 16'hFD42;    16'd61293: out <= 16'h0078;    16'd61294: out <= 16'h01E7;    16'd61295: out <= 16'h048B;
    16'd61296: out <= 16'h00E2;    16'd61297: out <= 16'h004F;    16'd61298: out <= 16'hFF54;    16'd61299: out <= 16'hFFA1;
    16'd61300: out <= 16'h071A;    16'd61301: out <= 16'hFE36;    16'd61302: out <= 16'h02D3;    16'd61303: out <= 16'hFCD8;
    16'd61304: out <= 16'h0321;    16'd61305: out <= 16'h01B2;    16'd61306: out <= 16'hFC65;    16'd61307: out <= 16'hFC8E;
    16'd61308: out <= 16'h0175;    16'd61309: out <= 16'h022A;    16'd61310: out <= 16'hF929;    16'd61311: out <= 16'h0698;
    16'd61312: out <= 16'h0803;    16'd61313: out <= 16'h01ED;    16'd61314: out <= 16'hFE9B;    16'd61315: out <= 16'hFCB8;
    16'd61316: out <= 16'hFE18;    16'd61317: out <= 16'h07CA;    16'd61318: out <= 16'h0008;    16'd61319: out <= 16'hFCA5;
    16'd61320: out <= 16'h03AA;    16'd61321: out <= 16'hFE50;    16'd61322: out <= 16'hF8CF;    16'd61323: out <= 16'h01A0;
    16'd61324: out <= 16'hFFA1;    16'd61325: out <= 16'h011F;    16'd61326: out <= 16'hFCBC;    16'd61327: out <= 16'hFB56;
    16'd61328: out <= 16'hFAF5;    16'd61329: out <= 16'h0342;    16'd61330: out <= 16'hFEBB;    16'd61331: out <= 16'hFA08;
    16'd61332: out <= 16'h015D;    16'd61333: out <= 16'h0082;    16'd61334: out <= 16'h052B;    16'd61335: out <= 16'hFF2D;
    16'd61336: out <= 16'h0708;    16'd61337: out <= 16'h05B7;    16'd61338: out <= 16'hFAE4;    16'd61339: out <= 16'hFDAE;
    16'd61340: out <= 16'hFF39;    16'd61341: out <= 16'h0222;    16'd61342: out <= 16'h009A;    16'd61343: out <= 16'hFE48;
    16'd61344: out <= 16'h012B;    16'd61345: out <= 16'h010B;    16'd61346: out <= 16'h0311;    16'd61347: out <= 16'hFCAF;
    16'd61348: out <= 16'h0142;    16'd61349: out <= 16'h081F;    16'd61350: out <= 16'hFEBA;    16'd61351: out <= 16'hF500;
    16'd61352: out <= 16'hFDA9;    16'd61353: out <= 16'hFD5B;    16'd61354: out <= 16'h0497;    16'd61355: out <= 16'h0140;
    16'd61356: out <= 16'h0656;    16'd61357: out <= 16'h055C;    16'd61358: out <= 16'h097A;    16'd61359: out <= 16'h039D;
    16'd61360: out <= 16'h0616;    16'd61361: out <= 16'h07B1;    16'd61362: out <= 16'hFF7C;    16'd61363: out <= 16'h051A;
    16'd61364: out <= 16'h03EB;    16'd61365: out <= 16'h02B0;    16'd61366: out <= 16'h00C8;    16'd61367: out <= 16'h0642;
    16'd61368: out <= 16'h092F;    16'd61369: out <= 16'h032F;    16'd61370: out <= 16'hFFE6;    16'd61371: out <= 16'h0428;
    16'd61372: out <= 16'hFF69;    16'd61373: out <= 16'h0648;    16'd61374: out <= 16'h043E;    16'd61375: out <= 16'h0908;
    16'd61376: out <= 16'h032B;    16'd61377: out <= 16'h09CC;    16'd61378: out <= 16'h035C;    16'd61379: out <= 16'h03B1;
    16'd61380: out <= 16'h056C;    16'd61381: out <= 16'h0333;    16'd61382: out <= 16'hFD14;    16'd61383: out <= 16'h04F9;
    16'd61384: out <= 16'hFECB;    16'd61385: out <= 16'h050B;    16'd61386: out <= 16'hFFEC;    16'd61387: out <= 16'hFEC5;
    16'd61388: out <= 16'hFA9E;    16'd61389: out <= 16'h009E;    16'd61390: out <= 16'h0239;    16'd61391: out <= 16'hFD50;
    16'd61392: out <= 16'hFD23;    16'd61393: out <= 16'h004A;    16'd61394: out <= 16'h0000;    16'd61395: out <= 16'h0168;
    16'd61396: out <= 16'h0092;    16'd61397: out <= 16'h0313;    16'd61398: out <= 16'h009A;    16'd61399: out <= 16'h0362;
    16'd61400: out <= 16'hFC18;    16'd61401: out <= 16'hFD21;    16'd61402: out <= 16'hF96F;    16'd61403: out <= 16'hFCA9;
    16'd61404: out <= 16'h0209;    16'd61405: out <= 16'hFF48;    16'd61406: out <= 16'h04F6;    16'd61407: out <= 16'h00E0;
    16'd61408: out <= 16'hFFBA;    16'd61409: out <= 16'h028F;    16'd61410: out <= 16'h0180;    16'd61411: out <= 16'h002D;
    16'd61412: out <= 16'h033E;    16'd61413: out <= 16'hF895;    16'd61414: out <= 16'h0247;    16'd61415: out <= 16'h0419;
    16'd61416: out <= 16'hFBD0;    16'd61417: out <= 16'h0195;    16'd61418: out <= 16'hFD77;    16'd61419: out <= 16'h0037;
    16'd61420: out <= 16'hFFA9;    16'd61421: out <= 16'h078D;    16'd61422: out <= 16'hFF8A;    16'd61423: out <= 16'hFF8B;
    16'd61424: out <= 16'hFA79;    16'd61425: out <= 16'h0215;    16'd61426: out <= 16'h095A;    16'd61427: out <= 16'hFE92;
    16'd61428: out <= 16'hFBE3;    16'd61429: out <= 16'h0479;    16'd61430: out <= 16'h01CA;    16'd61431: out <= 16'h016E;
    16'd61432: out <= 16'hFE02;    16'd61433: out <= 16'h03E1;    16'd61434: out <= 16'h00A1;    16'd61435: out <= 16'hFDA8;
    16'd61436: out <= 16'hFB35;    16'd61437: out <= 16'h001E;    16'd61438: out <= 16'hFB3F;    16'd61439: out <= 16'h086A;
    16'd61440: out <= 16'h06CC;    16'd61441: out <= 16'hF7CC;    16'd61442: out <= 16'h01B3;    16'd61443: out <= 16'hF9E7;
    16'd61444: out <= 16'hFE79;    16'd61445: out <= 16'hFD28;    16'd61446: out <= 16'hFDEE;    16'd61447: out <= 16'h02AB;
    16'd61448: out <= 16'h0767;    16'd61449: out <= 16'hFB83;    16'd61450: out <= 16'h0135;    16'd61451: out <= 16'hFD55;
    16'd61452: out <= 16'hFCED;    16'd61453: out <= 16'hFCEB;    16'd61454: out <= 16'hF9B0;    16'd61455: out <= 16'h0086;
    16'd61456: out <= 16'h0225;    16'd61457: out <= 16'h02A1;    16'd61458: out <= 16'h018C;    16'd61459: out <= 16'hFC1A;
    16'd61460: out <= 16'hFB84;    16'd61461: out <= 16'hFC41;    16'd61462: out <= 16'h015A;    16'd61463: out <= 16'h0404;
    16'd61464: out <= 16'h07A1;    16'd61465: out <= 16'hFF34;    16'd61466: out <= 16'h0418;    16'd61467: out <= 16'hFE41;
    16'd61468: out <= 16'h0225;    16'd61469: out <= 16'hFF9B;    16'd61470: out <= 16'h0005;    16'd61471: out <= 16'hF952;
    16'd61472: out <= 16'h00EB;    16'd61473: out <= 16'h0211;    16'd61474: out <= 16'h0676;    16'd61475: out <= 16'hFF20;
    16'd61476: out <= 16'h0261;    16'd61477: out <= 16'h0003;    16'd61478: out <= 16'hFF0F;    16'd61479: out <= 16'hFB4B;
    16'd61480: out <= 16'hFF5A;    16'd61481: out <= 16'hFD5A;    16'd61482: out <= 16'hF981;    16'd61483: out <= 16'hFAAF;
    16'd61484: out <= 16'h00CB;    16'd61485: out <= 16'h06FE;    16'd61486: out <= 16'h0795;    16'd61487: out <= 16'h04CE;
    16'd61488: out <= 16'h07BF;    16'd61489: out <= 16'h0587;    16'd61490: out <= 16'h00C1;    16'd61491: out <= 16'h107B;
    16'd61492: out <= 16'h02F1;    16'd61493: out <= 16'h0350;    16'd61494: out <= 16'hFCC8;    16'd61495: out <= 16'h01D5;
    16'd61496: out <= 16'h0104;    16'd61497: out <= 16'h049E;    16'd61498: out <= 16'h008C;    16'd61499: out <= 16'h0567;
    16'd61500: out <= 16'h09A6;    16'd61501: out <= 16'h029D;    16'd61502: out <= 16'h082C;    16'd61503: out <= 16'h001D;
    16'd61504: out <= 16'h0372;    16'd61505: out <= 16'h0A41;    16'd61506: out <= 16'h017E;    16'd61507: out <= 16'hFCF7;
    16'd61508: out <= 16'h08AB;    16'd61509: out <= 16'h0149;    16'd61510: out <= 16'hFEFA;    16'd61511: out <= 16'hFD2C;
    16'd61512: out <= 16'h04F8;    16'd61513: out <= 16'h0308;    16'd61514: out <= 16'h09EE;    16'd61515: out <= 16'h08EB;
    16'd61516: out <= 16'h0308;    16'd61517: out <= 16'h049E;    16'd61518: out <= 16'h06D7;    16'd61519: out <= 16'h03D8;
    16'd61520: out <= 16'hF81C;    16'd61521: out <= 16'h0620;    16'd61522: out <= 16'hFF7E;    16'd61523: out <= 16'hFE8D;
    16'd61524: out <= 16'hFFE0;    16'd61525: out <= 16'hFD9D;    16'd61526: out <= 16'hFE52;    16'd61527: out <= 16'h02E1;
    16'd61528: out <= 16'hFB57;    16'd61529: out <= 16'hFBF8;    16'd61530: out <= 16'h004A;    16'd61531: out <= 16'hFE95;
    16'd61532: out <= 16'hFF92;    16'd61533: out <= 16'h027E;    16'd61534: out <= 16'hFF52;    16'd61535: out <= 16'h089D;
    16'd61536: out <= 16'h009D;    16'd61537: out <= 16'hFDC1;    16'd61538: out <= 16'hFBC3;    16'd61539: out <= 16'h01EF;
    16'd61540: out <= 16'h0626;    16'd61541: out <= 16'h0411;    16'd61542: out <= 16'hF6D2;    16'd61543: out <= 16'h03A3;
    16'd61544: out <= 16'hF732;    16'd61545: out <= 16'hF64F;    16'd61546: out <= 16'h0274;    16'd61547: out <= 16'hFED4;
    16'd61548: out <= 16'h009D;    16'd61549: out <= 16'hFF7F;    16'd61550: out <= 16'h031C;    16'd61551: out <= 16'hFD44;
    16'd61552: out <= 16'h04AA;    16'd61553: out <= 16'h00C7;    16'd61554: out <= 16'h0371;    16'd61555: out <= 16'h01FB;
    16'd61556: out <= 16'hF83D;    16'd61557: out <= 16'h060D;    16'd61558: out <= 16'hFDB1;    16'd61559: out <= 16'hFF6D;
    16'd61560: out <= 16'hF93B;    16'd61561: out <= 16'h03A0;    16'd61562: out <= 16'h042C;    16'd61563: out <= 16'hFDA0;
    16'd61564: out <= 16'hFF4F;    16'd61565: out <= 16'hFE35;    16'd61566: out <= 16'h077C;    16'd61567: out <= 16'hFE6E;
    16'd61568: out <= 16'hFEBD;    16'd61569: out <= 16'h04BA;    16'd61570: out <= 16'h0034;    16'd61571: out <= 16'hF9EF;
    16'd61572: out <= 16'h005F;    16'd61573: out <= 16'h0226;    16'd61574: out <= 16'hFC18;    16'd61575: out <= 16'hF5AD;
    16'd61576: out <= 16'h00C9;    16'd61577: out <= 16'hFAF4;    16'd61578: out <= 16'hFF3B;    16'd61579: out <= 16'hFC8C;
    16'd61580: out <= 16'hFED9;    16'd61581: out <= 16'h04E6;    16'd61582: out <= 16'h0003;    16'd61583: out <= 16'h02AD;
    16'd61584: out <= 16'h05B4;    16'd61585: out <= 16'h0486;    16'd61586: out <= 16'hFFDC;    16'd61587: out <= 16'h03AA;
    16'd61588: out <= 16'hFBA5;    16'd61589: out <= 16'h0335;    16'd61590: out <= 16'h0199;    16'd61591: out <= 16'hFA95;
    16'd61592: out <= 16'hF5DE;    16'd61593: out <= 16'hFE72;    16'd61594: out <= 16'h0465;    16'd61595: out <= 16'hFF70;
    16'd61596: out <= 16'hF9FD;    16'd61597: out <= 16'hF996;    16'd61598: out <= 16'h01D2;    16'd61599: out <= 16'hFF6A;
    16'd61600: out <= 16'h0089;    16'd61601: out <= 16'h007D;    16'd61602: out <= 16'h00B5;    16'd61603: out <= 16'hFEB8;
    16'd61604: out <= 16'hFB4B;    16'd61605: out <= 16'hFD18;    16'd61606: out <= 16'hFFE1;    16'd61607: out <= 16'h062A;
    16'd61608: out <= 16'h0035;    16'd61609: out <= 16'h0161;    16'd61610: out <= 16'h06A9;    16'd61611: out <= 16'h008C;
    16'd61612: out <= 16'hFFAB;    16'd61613: out <= 16'h001F;    16'd61614: out <= 16'h04E1;    16'd61615: out <= 16'h064B;
    16'd61616: out <= 16'hFE25;    16'd61617: out <= 16'h011D;    16'd61618: out <= 16'h087A;    16'd61619: out <= 16'h032A;
    16'd61620: out <= 16'h063A;    16'd61621: out <= 16'hFFF4;    16'd61622: out <= 16'h0373;    16'd61623: out <= 16'h0333;
    16'd61624: out <= 16'h036A;    16'd61625: out <= 16'hFDC3;    16'd61626: out <= 16'h008D;    16'd61627: out <= 16'hFF1D;
    16'd61628: out <= 16'h0446;    16'd61629: out <= 16'h052B;    16'd61630: out <= 16'h099A;    16'd61631: out <= 16'h03D5;
    16'd61632: out <= 16'h0603;    16'd61633: out <= 16'h05F0;    16'd61634: out <= 16'h04EC;    16'd61635: out <= 16'h0825;
    16'd61636: out <= 16'h08BA;    16'd61637: out <= 16'h03A2;    16'd61638: out <= 16'h03C5;    16'd61639: out <= 16'h0615;
    16'd61640: out <= 16'hFEE8;    16'd61641: out <= 16'hFDB7;    16'd61642: out <= 16'hFC3A;    16'd61643: out <= 16'h0538;
    16'd61644: out <= 16'h035A;    16'd61645: out <= 16'h0141;    16'd61646: out <= 16'hFE66;    16'd61647: out <= 16'h0271;
    16'd61648: out <= 16'h0130;    16'd61649: out <= 16'hF9E3;    16'd61650: out <= 16'h0324;    16'd61651: out <= 16'h0A84;
    16'd61652: out <= 16'h0002;    16'd61653: out <= 16'h057A;    16'd61654: out <= 16'hFD81;    16'd61655: out <= 16'h08B8;
    16'd61656: out <= 16'h024D;    16'd61657: out <= 16'h012A;    16'd61658: out <= 16'h056F;    16'd61659: out <= 16'hFE44;
    16'd61660: out <= 16'h0262;    16'd61661: out <= 16'h0532;    16'd61662: out <= 16'hFEA7;    16'd61663: out <= 16'hF9A7;
    16'd61664: out <= 16'hFD0A;    16'd61665: out <= 16'hFE16;    16'd61666: out <= 16'h03F8;    16'd61667: out <= 16'hFA19;
    16'd61668: out <= 16'h017E;    16'd61669: out <= 16'h06F2;    16'd61670: out <= 16'h017B;    16'd61671: out <= 16'hFE7B;
    16'd61672: out <= 16'hFF27;    16'd61673: out <= 16'hF61D;    16'd61674: out <= 16'h0343;    16'd61675: out <= 16'hFD86;
    16'd61676: out <= 16'hFCC0;    16'd61677: out <= 16'h0150;    16'd61678: out <= 16'h0056;    16'd61679: out <= 16'hFDA2;
    16'd61680: out <= 16'h03AB;    16'd61681: out <= 16'h0209;    16'd61682: out <= 16'hF702;    16'd61683: out <= 16'h0036;
    16'd61684: out <= 16'hFE88;    16'd61685: out <= 16'hFFA0;    16'd61686: out <= 16'hFDC6;    16'd61687: out <= 16'hFD7C;
    16'd61688: out <= 16'h0639;    16'd61689: out <= 16'hFE8E;    16'd61690: out <= 16'hFA69;    16'd61691: out <= 16'h0108;
    16'd61692: out <= 16'hFC43;    16'd61693: out <= 16'hFB3D;    16'd61694: out <= 16'h015B;    16'd61695: out <= 16'hFE1B;
    16'd61696: out <= 16'hFE91;    16'd61697: out <= 16'hFE4E;    16'd61698: out <= 16'hFD6D;    16'd61699: out <= 16'h0128;
    16'd61700: out <= 16'hFFF8;    16'd61701: out <= 16'hFA3F;    16'd61702: out <= 16'h04D1;    16'd61703: out <= 16'hFE74;
    16'd61704: out <= 16'hFC84;    16'd61705: out <= 16'hFF46;    16'd61706: out <= 16'hFFCE;    16'd61707: out <= 16'h0626;
    16'd61708: out <= 16'h0462;    16'd61709: out <= 16'h056B;    16'd61710: out <= 16'hFEAC;    16'd61711: out <= 16'hFEE7;
    16'd61712: out <= 16'h0385;    16'd61713: out <= 16'h0080;    16'd61714: out <= 16'hFC2F;    16'd61715: out <= 16'hF9E3;
    16'd61716: out <= 16'hF8DC;    16'd61717: out <= 16'h079C;    16'd61718: out <= 16'hF955;    16'd61719: out <= 16'h021C;
    16'd61720: out <= 16'h04D9;    16'd61721: out <= 16'h01CE;    16'd61722: out <= 16'hFF3C;    16'd61723: out <= 16'hFEDA;
    16'd61724: out <= 16'h057B;    16'd61725: out <= 16'hFB45;    16'd61726: out <= 16'h030C;    16'd61727: out <= 16'h0139;
    16'd61728: out <= 16'hFD2F;    16'd61729: out <= 16'h010A;    16'd61730: out <= 16'h0428;    16'd61731: out <= 16'h0470;
    16'd61732: out <= 16'h02E7;    16'd61733: out <= 16'h073D;    16'd61734: out <= 16'h01CB;    16'd61735: out <= 16'hFC39;
    16'd61736: out <= 16'hFEA2;    16'd61737: out <= 16'h03E2;    16'd61738: out <= 16'hFFA4;    16'd61739: out <= 16'hFE5C;
    16'd61740: out <= 16'hFC63;    16'd61741: out <= 16'h0693;    16'd61742: out <= 16'h0068;    16'd61743: out <= 16'h0514;
    16'd61744: out <= 16'h048D;    16'd61745: out <= 16'h0173;    16'd61746: out <= 16'h0A72;    16'd61747: out <= 16'h0743;
    16'd61748: out <= 16'h0696;    16'd61749: out <= 16'h031D;    16'd61750: out <= 16'h0834;    16'd61751: out <= 16'hFF0F;
    16'd61752: out <= 16'h02A1;    16'd61753: out <= 16'h03FD;    16'd61754: out <= 16'h048A;    16'd61755: out <= 16'h0434;
    16'd61756: out <= 16'h0547;    16'd61757: out <= 16'h08F7;    16'd61758: out <= 16'h0672;    16'd61759: out <= 16'h05F6;
    16'd61760: out <= 16'hFEB4;    16'd61761: out <= 16'h067D;    16'd61762: out <= 16'h0649;    16'd61763: out <= 16'h098D;
    16'd61764: out <= 16'h0AE7;    16'd61765: out <= 16'hFFDA;    16'd61766: out <= 16'h048C;    16'd61767: out <= 16'h0818;
    16'd61768: out <= 16'h01D6;    16'd61769: out <= 16'hFF4B;    16'd61770: out <= 16'hFC2A;    16'd61771: out <= 16'h03B5;
    16'd61772: out <= 16'hFCEA;    16'd61773: out <= 16'h01A1;    16'd61774: out <= 16'hFEF5;    16'd61775: out <= 16'h0456;
    16'd61776: out <= 16'hFB4D;    16'd61777: out <= 16'h017A;    16'd61778: out <= 16'h0223;    16'd61779: out <= 16'hFCD7;
    16'd61780: out <= 16'hF7A2;    16'd61781: out <= 16'h0185;    16'd61782: out <= 16'h009A;    16'd61783: out <= 16'hFEB0;
    16'd61784: out <= 16'hFC5E;    16'd61785: out <= 16'h0206;    16'd61786: out <= 16'hFFA7;    16'd61787: out <= 16'hFFBD;
    16'd61788: out <= 16'h01D5;    16'd61789: out <= 16'h05C7;    16'd61790: out <= 16'h000B;    16'd61791: out <= 16'hFE86;
    16'd61792: out <= 16'h02F0;    16'd61793: out <= 16'hFBC9;    16'd61794: out <= 16'h00F1;    16'd61795: out <= 16'hFB43;
    16'd61796: out <= 16'hF6DE;    16'd61797: out <= 16'hFD2E;    16'd61798: out <= 16'hFFC1;    16'd61799: out <= 16'hFA54;
    16'd61800: out <= 16'h0336;    16'd61801: out <= 16'h0188;    16'd61802: out <= 16'hFD68;    16'd61803: out <= 16'hFDE2;
    16'd61804: out <= 16'h003B;    16'd61805: out <= 16'h01E5;    16'd61806: out <= 16'hFE30;    16'd61807: out <= 16'hFDDC;
    16'd61808: out <= 16'hF468;    16'd61809: out <= 16'hF9A6;    16'd61810: out <= 16'hFAEE;    16'd61811: out <= 16'hFD33;
    16'd61812: out <= 16'h0397;    16'd61813: out <= 16'h0446;    16'd61814: out <= 16'h0332;    16'd61815: out <= 16'hFFD2;
    16'd61816: out <= 16'hF887;    16'd61817: out <= 16'hFD2D;    16'd61818: out <= 16'hFAD4;    16'd61819: out <= 16'h0554;
    16'd61820: out <= 16'h0112;    16'd61821: out <= 16'h0578;    16'd61822: out <= 16'h0090;    16'd61823: out <= 16'hFB3D;
    16'd61824: out <= 16'h01C1;    16'd61825: out <= 16'h0370;    16'd61826: out <= 16'hFECE;    16'd61827: out <= 16'hFF02;
    16'd61828: out <= 16'h0588;    16'd61829: out <= 16'h00D7;    16'd61830: out <= 16'h01D8;    16'd61831: out <= 16'hFB2D;
    16'd61832: out <= 16'h084F;    16'd61833: out <= 16'hFF51;    16'd61834: out <= 16'h0255;    16'd61835: out <= 16'hFB84;
    16'd61836: out <= 16'hFED6;    16'd61837: out <= 16'h04E2;    16'd61838: out <= 16'h05B0;    16'd61839: out <= 16'hFEB3;
    16'd61840: out <= 16'hFEED;    16'd61841: out <= 16'hF9FD;    16'd61842: out <= 16'h010F;    16'd61843: out <= 16'hFEE8;
    16'd61844: out <= 16'h0151;    16'd61845: out <= 16'hFE89;    16'd61846: out <= 16'hFD4B;    16'd61847: out <= 16'h04B1;
    16'd61848: out <= 16'hFDA2;    16'd61849: out <= 16'h028C;    16'd61850: out <= 16'h0256;    16'd61851: out <= 16'hFFA0;
    16'd61852: out <= 16'hFB46;    16'd61853: out <= 16'hFF30;    16'd61854: out <= 16'h02FD;    16'd61855: out <= 16'h03F7;
    16'd61856: out <= 16'h027C;    16'd61857: out <= 16'h02C5;    16'd61858: out <= 16'h02FD;    16'd61859: out <= 16'hF977;
    16'd61860: out <= 16'hFF03;    16'd61861: out <= 16'h07A1;    16'd61862: out <= 16'h083A;    16'd61863: out <= 16'h00E1;
    16'd61864: out <= 16'hFCCB;    16'd61865: out <= 16'h07A0;    16'd61866: out <= 16'h07A6;    16'd61867: out <= 16'hFF4E;
    16'd61868: out <= 16'h0AEE;    16'd61869: out <= 16'hFC14;    16'd61870: out <= 16'h02B9;    16'd61871: out <= 16'h0308;
    16'd61872: out <= 16'h0232;    16'd61873: out <= 16'h0778;    16'd61874: out <= 16'h0240;    16'd61875: out <= 16'h004B;
    16'd61876: out <= 16'h0331;    16'd61877: out <= 16'h0500;    16'd61878: out <= 16'hFFE2;    16'd61879: out <= 16'h0D99;
    16'd61880: out <= 16'hFD7C;    16'd61881: out <= 16'h0415;    16'd61882: out <= 16'h099A;    16'd61883: out <= 16'h0732;
    16'd61884: out <= 16'h0055;    16'd61885: out <= 16'h08E8;    16'd61886: out <= 16'h0495;    16'd61887: out <= 16'h0359;
    16'd61888: out <= 16'h054D;    16'd61889: out <= 16'hFEFC;    16'd61890: out <= 16'h0819;    16'd61891: out <= 16'h0BB8;
    16'd61892: out <= 16'h0176;    16'd61893: out <= 16'h0312;    16'd61894: out <= 16'hFE17;    16'd61895: out <= 16'h00B6;
    16'd61896: out <= 16'hFFA7;    16'd61897: out <= 16'h00A9;    16'd61898: out <= 16'h03C4;    16'd61899: out <= 16'h030A;
    16'd61900: out <= 16'h0317;    16'd61901: out <= 16'h030F;    16'd61902: out <= 16'hFD4D;    16'd61903: out <= 16'hFB9B;
    16'd61904: out <= 16'h021A;    16'd61905: out <= 16'hFE3E;    16'd61906: out <= 16'h081D;    16'd61907: out <= 16'h0011;
    16'd61908: out <= 16'hFE8A;    16'd61909: out <= 16'h015B;    16'd61910: out <= 16'hFDB6;    16'd61911: out <= 16'h0049;
    16'd61912: out <= 16'h015E;    16'd61913: out <= 16'hFC24;    16'd61914: out <= 16'h0266;    16'd61915: out <= 16'h069B;
    16'd61916: out <= 16'hFABA;    16'd61917: out <= 16'h02C5;    16'd61918: out <= 16'h00DA;    16'd61919: out <= 16'h0074;
    16'd61920: out <= 16'h0372;    16'd61921: out <= 16'h0681;    16'd61922: out <= 16'hFCDA;    16'd61923: out <= 16'h0083;
    16'd61924: out <= 16'hFCC0;    16'd61925: out <= 16'hFD2B;    16'd61926: out <= 16'hFCDB;    16'd61927: out <= 16'hFC65;
    16'd61928: out <= 16'hFCA3;    16'd61929: out <= 16'hFF82;    16'd61930: out <= 16'h02F8;    16'd61931: out <= 16'hFE09;
    16'd61932: out <= 16'h02EE;    16'd61933: out <= 16'h00DA;    16'd61934: out <= 16'hFE71;    16'd61935: out <= 16'h03EA;
    16'd61936: out <= 16'h03D2;    16'd61937: out <= 16'h045A;    16'd61938: out <= 16'h0899;    16'd61939: out <= 16'h03CD;
    16'd61940: out <= 16'h007C;    16'd61941: out <= 16'h022E;    16'd61942: out <= 16'h01D2;    16'd61943: out <= 16'h018D;
    16'd61944: out <= 16'hFFD2;    16'd61945: out <= 16'h000B;    16'd61946: out <= 16'h0601;    16'd61947: out <= 16'hFB9A;
    16'd61948: out <= 16'hF912;    16'd61949: out <= 16'hFC4B;    16'd61950: out <= 16'h0429;    16'd61951: out <= 16'h0335;
    16'd61952: out <= 16'hFD07;    16'd61953: out <= 16'h039C;    16'd61954: out <= 16'h0040;    16'd61955: out <= 16'hFFC2;
    16'd61956: out <= 16'hFFBD;    16'd61957: out <= 16'hFDEB;    16'd61958: out <= 16'h043A;    16'd61959: out <= 16'h029E;
    16'd61960: out <= 16'hFE9D;    16'd61961: out <= 16'hFDB3;    16'd61962: out <= 16'hFE89;    16'd61963: out <= 16'hFD58;
    16'd61964: out <= 16'hF893;    16'd61965: out <= 16'hFD91;    16'd61966: out <= 16'h04E1;    16'd61967: out <= 16'hFF89;
    16'd61968: out <= 16'h0047;    16'd61969: out <= 16'hFCCB;    16'd61970: out <= 16'hFEA4;    16'd61971: out <= 16'hF8B7;
    16'd61972: out <= 16'hFA08;    16'd61973: out <= 16'h023D;    16'd61974: out <= 16'hFD24;    16'd61975: out <= 16'h023A;
    16'd61976: out <= 16'hFC5C;    16'd61977: out <= 16'hFAB7;    16'd61978: out <= 16'hFFD7;    16'd61979: out <= 16'h00B2;
    16'd61980: out <= 16'hFE4F;    16'd61981: out <= 16'hF8C2;    16'd61982: out <= 16'h03C6;    16'd61983: out <= 16'hFFBF;
    16'd61984: out <= 16'hFC82;    16'd61985: out <= 16'h003F;    16'd61986: out <= 16'hFD8A;    16'd61987: out <= 16'h00EC;
    16'd61988: out <= 16'hFFC6;    16'd61989: out <= 16'hFB77;    16'd61990: out <= 16'h0414;    16'd61991: out <= 16'h0122;
    16'd61992: out <= 16'hFDF6;    16'd61993: out <= 16'hFEA6;    16'd61994: out <= 16'hFD8D;    16'd61995: out <= 16'h026F;
    16'd61996: out <= 16'hFCCD;    16'd61997: out <= 16'h0100;    16'd61998: out <= 16'h0CD8;    16'd61999: out <= 16'h0213;
    16'd62000: out <= 16'h06AE;    16'd62001: out <= 16'h06EF;    16'd62002: out <= 16'h04DD;    16'd62003: out <= 16'h0096;
    16'd62004: out <= 16'h05CA;    16'd62005: out <= 16'h022F;    16'd62006: out <= 16'hFC09;    16'd62007: out <= 16'h019D;
    16'd62008: out <= 16'h0920;    16'd62009: out <= 16'h00F4;    16'd62010: out <= 16'h061B;    16'd62011: out <= 16'h09E5;
    16'd62012: out <= 16'h052B;    16'd62013: out <= 16'h025F;    16'd62014: out <= 16'h0933;    16'd62015: out <= 16'h0A64;
    16'd62016: out <= 16'h001B;    16'd62017: out <= 16'h0257;    16'd62018: out <= 16'h091E;    16'd62019: out <= 16'h03B2;
    16'd62020: out <= 16'hFDF5;    16'd62021: out <= 16'hFE09;    16'd62022: out <= 16'h05DE;    16'd62023: out <= 16'hFE28;
    16'd62024: out <= 16'h03B4;    16'd62025: out <= 16'h0063;    16'd62026: out <= 16'hFD64;    16'd62027: out <= 16'hFDDC;
    16'd62028: out <= 16'h05E5;    16'd62029: out <= 16'h03E4;    16'd62030: out <= 16'h031A;    16'd62031: out <= 16'h0153;
    16'd62032: out <= 16'hFD56;    16'd62033: out <= 16'h071F;    16'd62034: out <= 16'h0237;    16'd62035: out <= 16'h044C;
    16'd62036: out <= 16'hF8B0;    16'd62037: out <= 16'h04CF;    16'd62038: out <= 16'hFB5A;    16'd62039: out <= 16'hFA37;
    16'd62040: out <= 16'hFB5E;    16'd62041: out <= 16'hF6F4;    16'd62042: out <= 16'h0342;    16'd62043: out <= 16'h01B3;
    16'd62044: out <= 16'hFC18;    16'd62045: out <= 16'hFFB9;    16'd62046: out <= 16'hFF1B;    16'd62047: out <= 16'h0429;
    16'd62048: out <= 16'hFA50;    16'd62049: out <= 16'h0221;    16'd62050: out <= 16'hFD95;    16'd62051: out <= 16'hFE6E;
    16'd62052: out <= 16'h00E8;    16'd62053: out <= 16'h04A6;    16'd62054: out <= 16'h00BE;    16'd62055: out <= 16'h015B;
    16'd62056: out <= 16'h0223;    16'd62057: out <= 16'h0290;    16'd62058: out <= 16'h0201;    16'd62059: out <= 16'hF7BF;
    16'd62060: out <= 16'h056C;    16'd62061: out <= 16'hFFBE;    16'd62062: out <= 16'hFA23;    16'd62063: out <= 16'h0182;
    16'd62064: out <= 16'hFEDE;    16'd62065: out <= 16'hF841;    16'd62066: out <= 16'h033E;    16'd62067: out <= 16'hFB3C;
    16'd62068: out <= 16'h00FD;    16'd62069: out <= 16'h0448;    16'd62070: out <= 16'h004E;    16'd62071: out <= 16'h0326;
    16'd62072: out <= 16'hFD9E;    16'd62073: out <= 16'h06CB;    16'd62074: out <= 16'hFF3F;    16'd62075: out <= 16'h0634;
    16'd62076: out <= 16'hFA5C;    16'd62077: out <= 16'hFDE0;    16'd62078: out <= 16'h062A;    16'd62079: out <= 16'hFABA;
    16'd62080: out <= 16'hFC3A;    16'd62081: out <= 16'hFD9A;    16'd62082: out <= 16'h0363;    16'd62083: out <= 16'h0503;
    16'd62084: out <= 16'h03CA;    16'd62085: out <= 16'h00E7;    16'd62086: out <= 16'h0319;    16'd62087: out <= 16'h07BA;
    16'd62088: out <= 16'hF7B6;    16'd62089: out <= 16'hFF54;    16'd62090: out <= 16'h0642;    16'd62091: out <= 16'hFB50;
    16'd62092: out <= 16'h03E0;    16'd62093: out <= 16'hFD19;    16'd62094: out <= 16'hF889;    16'd62095: out <= 16'hFBAE;
    16'd62096: out <= 16'hFCE7;    16'd62097: out <= 16'h012B;    16'd62098: out <= 16'hFB04;    16'd62099: out <= 16'hFAB3;
    16'd62100: out <= 16'h0092;    16'd62101: out <= 16'hFE56;    16'd62102: out <= 16'hFE03;    16'd62103: out <= 16'h06C6;
    16'd62104: out <= 16'hF916;    16'd62105: out <= 16'h0143;    16'd62106: out <= 16'hF983;    16'd62107: out <= 16'hFDF2;
    16'd62108: out <= 16'h0009;    16'd62109: out <= 16'hFF25;    16'd62110: out <= 16'hFDB0;    16'd62111: out <= 16'h06B8;
    16'd62112: out <= 16'hFAE0;    16'd62113: out <= 16'hFB4F;    16'd62114: out <= 16'hFEEA;    16'd62115: out <= 16'hFF30;
    16'd62116: out <= 16'h0208;    16'd62117: out <= 16'hFD3B;    16'd62118: out <= 16'h011B;    16'd62119: out <= 16'hFADD;
    16'd62120: out <= 16'hF987;    16'd62121: out <= 16'h0252;    16'd62122: out <= 16'h0221;    16'd62123: out <= 16'h0615;
    16'd62124: out <= 16'h0361;    16'd62125: out <= 16'h064B;    16'd62126: out <= 16'h01A2;    16'd62127: out <= 16'h0135;
    16'd62128: out <= 16'h0160;    16'd62129: out <= 16'h08A2;    16'd62130: out <= 16'h0313;    16'd62131: out <= 16'hFC3F;
    16'd62132: out <= 16'h03F4;    16'd62133: out <= 16'h0A52;    16'd62134: out <= 16'h0519;    16'd62135: out <= 16'h0997;
    16'd62136: out <= 16'h06BB;    16'd62137: out <= 16'hFBBA;    16'd62138: out <= 16'h0337;    16'd62139: out <= 16'h0518;
    16'd62140: out <= 16'h0246;    16'd62141: out <= 16'h0562;    16'd62142: out <= 16'h00CE;    16'd62143: out <= 16'h0165;
    16'd62144: out <= 16'h09C6;    16'd62145: out <= 16'h0814;    16'd62146: out <= 16'h06D4;    16'd62147: out <= 16'hFE77;
    16'd62148: out <= 16'hFF3A;    16'd62149: out <= 16'hFD95;    16'd62150: out <= 16'hFE03;    16'd62151: out <= 16'hFC09;
    16'd62152: out <= 16'h00F6;    16'd62153: out <= 16'h0A48;    16'd62154: out <= 16'hF901;    16'd62155: out <= 16'hFC4A;
    16'd62156: out <= 16'h05E0;    16'd62157: out <= 16'h0244;    16'd62158: out <= 16'h0434;    16'd62159: out <= 16'hF7CF;
    16'd62160: out <= 16'h0186;    16'd62161: out <= 16'h0029;    16'd62162: out <= 16'hFD89;    16'd62163: out <= 16'h004A;
    16'd62164: out <= 16'hFFAA;    16'd62165: out <= 16'hFF20;    16'd62166: out <= 16'hFA35;    16'd62167: out <= 16'h0415;
    16'd62168: out <= 16'h026A;    16'd62169: out <= 16'h0391;    16'd62170: out <= 16'h078A;    16'd62171: out <= 16'h0470;
    16'd62172: out <= 16'hFD89;    16'd62173: out <= 16'hF97E;    16'd62174: out <= 16'hFF93;    16'd62175: out <= 16'hFFDF;
    16'd62176: out <= 16'h05B0;    16'd62177: out <= 16'hFECA;    16'd62178: out <= 16'hFCEA;    16'd62179: out <= 16'hFA44;
    16'd62180: out <= 16'h0344;    16'd62181: out <= 16'hFB98;    16'd62182: out <= 16'h03B7;    16'd62183: out <= 16'hF76D;
    16'd62184: out <= 16'h005B;    16'd62185: out <= 16'hFFDB;    16'd62186: out <= 16'hFF04;    16'd62187: out <= 16'h002E;
    16'd62188: out <= 16'h0752;    16'd62189: out <= 16'h036C;    16'd62190: out <= 16'h03BF;    16'd62191: out <= 16'hFFAA;
    16'd62192: out <= 16'hFD99;    16'd62193: out <= 16'hFB70;    16'd62194: out <= 16'h042F;    16'd62195: out <= 16'h03F0;
    16'd62196: out <= 16'hFBCB;    16'd62197: out <= 16'hFE8B;    16'd62198: out <= 16'hFD43;    16'd62199: out <= 16'h0822;
    16'd62200: out <= 16'h0061;    16'd62201: out <= 16'h08A1;    16'd62202: out <= 16'h033C;    16'd62203: out <= 16'h00E9;
    16'd62204: out <= 16'h0565;    16'd62205: out <= 16'hFCAB;    16'd62206: out <= 16'hF88B;    16'd62207: out <= 16'h0324;
    16'd62208: out <= 16'h01EE;    16'd62209: out <= 16'h0388;    16'd62210: out <= 16'h03E1;    16'd62211: out <= 16'h05D4;
    16'd62212: out <= 16'hFA81;    16'd62213: out <= 16'hFBCD;    16'd62214: out <= 16'h0587;    16'd62215: out <= 16'hFEC6;
    16'd62216: out <= 16'hFE58;    16'd62217: out <= 16'hFF7F;    16'd62218: out <= 16'hF95D;    16'd62219: out <= 16'h0349;
    16'd62220: out <= 16'hF9C2;    16'd62221: out <= 16'h0625;    16'd62222: out <= 16'hFE73;    16'd62223: out <= 16'hFE6A;
    16'd62224: out <= 16'hF8F4;    16'd62225: out <= 16'h0745;    16'd62226: out <= 16'h0254;    16'd62227: out <= 16'hFC1B;
    16'd62228: out <= 16'hFEAC;    16'd62229: out <= 16'h0013;    16'd62230: out <= 16'h03A3;    16'd62231: out <= 16'h00C4;
    16'd62232: out <= 16'h0533;    16'd62233: out <= 16'hF6CD;    16'd62234: out <= 16'h07FB;    16'd62235: out <= 16'h0027;
    16'd62236: out <= 16'hFCAB;    16'd62237: out <= 16'h04B6;    16'd62238: out <= 16'hFB31;    16'd62239: out <= 16'hFE66;
    16'd62240: out <= 16'h014E;    16'd62241: out <= 16'h0154;    16'd62242: out <= 16'hF67F;    16'd62243: out <= 16'h032E;
    16'd62244: out <= 16'hFB70;    16'd62245: out <= 16'h00C7;    16'd62246: out <= 16'hFCAC;    16'd62247: out <= 16'h00E2;
    16'd62248: out <= 16'hFFAD;    16'd62249: out <= 16'h01CF;    16'd62250: out <= 16'h0567;    16'd62251: out <= 16'h0183;
    16'd62252: out <= 16'h090C;    16'd62253: out <= 16'h0327;    16'd62254: out <= 16'h03E1;    16'd62255: out <= 16'h026C;
    16'd62256: out <= 16'h03E2;    16'd62257: out <= 16'h050F;    16'd62258: out <= 16'h003A;    16'd62259: out <= 16'h0869;
    16'd62260: out <= 16'h041B;    16'd62261: out <= 16'h0B19;    16'd62262: out <= 16'h04FE;    16'd62263: out <= 16'h048A;
    16'd62264: out <= 16'h0658;    16'd62265: out <= 16'h0328;    16'd62266: out <= 16'h0401;    16'd62267: out <= 16'h04CF;
    16'd62268: out <= 16'h07B6;    16'd62269: out <= 16'h002D;    16'd62270: out <= 16'h00F1;    16'd62271: out <= 16'h035A;
    16'd62272: out <= 16'h0931;    16'd62273: out <= 16'h03EA;    16'd62274: out <= 16'h0B36;    16'd62275: out <= 16'hFA4F;
    16'd62276: out <= 16'h0750;    16'd62277: out <= 16'h0196;    16'd62278: out <= 16'hFECC;    16'd62279: out <= 16'h0715;
    16'd62280: out <= 16'h0525;    16'd62281: out <= 16'h07B5;    16'd62282: out <= 16'h0656;    16'd62283: out <= 16'hFD3A;
    16'd62284: out <= 16'h063F;    16'd62285: out <= 16'h047B;    16'd62286: out <= 16'h05C8;    16'd62287: out <= 16'hFF42;
    16'd62288: out <= 16'hFBB6;    16'd62289: out <= 16'hFB02;    16'd62290: out <= 16'h00E9;    16'd62291: out <= 16'h08BE;
    16'd62292: out <= 16'h0555;    16'd62293: out <= 16'h00B2;    16'd62294: out <= 16'hFD7F;    16'd62295: out <= 16'h02C8;
    16'd62296: out <= 16'h0462;    16'd62297: out <= 16'h00F9;    16'd62298: out <= 16'h04FE;    16'd62299: out <= 16'h0394;
    16'd62300: out <= 16'h0948;    16'd62301: out <= 16'hFFE6;    16'd62302: out <= 16'hFD05;    16'd62303: out <= 16'h041B;
    16'd62304: out <= 16'h0221;    16'd62305: out <= 16'hFE38;    16'd62306: out <= 16'hFBC3;    16'd62307: out <= 16'hFEA2;
    16'd62308: out <= 16'h0399;    16'd62309: out <= 16'hFDC9;    16'd62310: out <= 16'h0071;    16'd62311: out <= 16'h02C5;
    16'd62312: out <= 16'hFD6F;    16'd62313: out <= 16'hFC29;    16'd62314: out <= 16'h00FD;    16'd62315: out <= 16'hFDE3;
    16'd62316: out <= 16'hFFFB;    16'd62317: out <= 16'hFDA3;    16'd62318: out <= 16'hFF1C;    16'd62319: out <= 16'h02DF;
    16'd62320: out <= 16'h02D1;    16'd62321: out <= 16'h0412;    16'd62322: out <= 16'h0567;    16'd62323: out <= 16'hF6F6;
    16'd62324: out <= 16'h0542;    16'd62325: out <= 16'h02A8;    16'd62326: out <= 16'h01BF;    16'd62327: out <= 16'hF8D2;
    16'd62328: out <= 16'h04FC;    16'd62329: out <= 16'hFA63;    16'd62330: out <= 16'hFF1C;    16'd62331: out <= 16'h00C2;
    16'd62332: out <= 16'h019E;    16'd62333: out <= 16'h0571;    16'd62334: out <= 16'h000D;    16'd62335: out <= 16'h024D;
    16'd62336: out <= 16'h0015;    16'd62337: out <= 16'h07EB;    16'd62338: out <= 16'h01D0;    16'd62339: out <= 16'h0265;
    16'd62340: out <= 16'h0286;    16'd62341: out <= 16'hF919;    16'd62342: out <= 16'hF8A4;    16'd62343: out <= 16'hFA85;
    16'd62344: out <= 16'hFC0F;    16'd62345: out <= 16'h01C0;    16'd62346: out <= 16'h006A;    16'd62347: out <= 16'h01FA;
    16'd62348: out <= 16'h0164;    16'd62349: out <= 16'hFDFE;    16'd62350: out <= 16'hFD03;    16'd62351: out <= 16'h01D5;
    16'd62352: out <= 16'hFDB8;    16'd62353: out <= 16'h036B;    16'd62354: out <= 16'h066C;    16'd62355: out <= 16'h0019;
    16'd62356: out <= 16'hFB79;    16'd62357: out <= 16'h00A0;    16'd62358: out <= 16'h058B;    16'd62359: out <= 16'hFD97;
    16'd62360: out <= 16'h0328;    16'd62361: out <= 16'hFA99;    16'd62362: out <= 16'h01FC;    16'd62363: out <= 16'h06BC;
    16'd62364: out <= 16'h0283;    16'd62365: out <= 16'h074A;    16'd62366: out <= 16'hFD52;    16'd62367: out <= 16'h01E4;
    16'd62368: out <= 16'h0696;    16'd62369: out <= 16'h0576;    16'd62370: out <= 16'h066C;    16'd62371: out <= 16'hFFD5;
    16'd62372: out <= 16'h0186;    16'd62373: out <= 16'hFC08;    16'd62374: out <= 16'h01AF;    16'd62375: out <= 16'h09BC;
    16'd62376: out <= 16'hF9A9;    16'd62377: out <= 16'h06FC;    16'd62378: out <= 16'h0503;    16'd62379: out <= 16'h0562;
    16'd62380: out <= 16'h005A;    16'd62381: out <= 16'hF9B9;    16'd62382: out <= 16'hFD93;    16'd62383: out <= 16'h06B4;
    16'd62384: out <= 16'h0486;    16'd62385: out <= 16'h083A;    16'd62386: out <= 16'h041A;    16'd62387: out <= 16'hFFEF;
    16'd62388: out <= 16'h08D9;    16'd62389: out <= 16'h00B0;    16'd62390: out <= 16'h028C;    16'd62391: out <= 16'h02E4;
    16'd62392: out <= 16'h07ED;    16'd62393: out <= 16'h07C6;    16'd62394: out <= 16'h08FF;    16'd62395: out <= 16'h0448;
    16'd62396: out <= 16'h075C;    16'd62397: out <= 16'h0521;    16'd62398: out <= 16'h0403;    16'd62399: out <= 16'h0226;
    16'd62400: out <= 16'h0782;    16'd62401: out <= 16'h0A56;    16'd62402: out <= 16'h0919;    16'd62403: out <= 16'h0101;
    16'd62404: out <= 16'h00A1;    16'd62405: out <= 16'h0106;    16'd62406: out <= 16'h018B;    16'd62407: out <= 16'h040C;
    16'd62408: out <= 16'h00E1;    16'd62409: out <= 16'hFF56;    16'd62410: out <= 16'hF7F6;    16'd62411: out <= 16'hFEDB;
    16'd62412: out <= 16'hFE51;    16'd62413: out <= 16'h019A;    16'd62414: out <= 16'h0045;    16'd62415: out <= 16'h0082;
    16'd62416: out <= 16'hFD3C;    16'd62417: out <= 16'hFFEF;    16'd62418: out <= 16'h01EF;    16'd62419: out <= 16'hFCB7;
    16'd62420: out <= 16'hF8F8;    16'd62421: out <= 16'hF645;    16'd62422: out <= 16'h0147;    16'd62423: out <= 16'hF3CE;
    16'd62424: out <= 16'hFC09;    16'd62425: out <= 16'hFCD4;    16'd62426: out <= 16'h05E1;    16'd62427: out <= 16'h07AC;
    16'd62428: out <= 16'h0886;    16'd62429: out <= 16'h00D3;    16'd62430: out <= 16'hFCA9;    16'd62431: out <= 16'h01DA;
    16'd62432: out <= 16'h0293;    16'd62433: out <= 16'hFA00;    16'd62434: out <= 16'hFACF;    16'd62435: out <= 16'h0381;
    16'd62436: out <= 16'hFF37;    16'd62437: out <= 16'h03CC;    16'd62438: out <= 16'h0578;    16'd62439: out <= 16'h00A2;
    16'd62440: out <= 16'h0042;    16'd62441: out <= 16'hFFE9;    16'd62442: out <= 16'h0485;    16'd62443: out <= 16'h0831;
    16'd62444: out <= 16'h02B4;    16'd62445: out <= 16'hFE6F;    16'd62446: out <= 16'h03D0;    16'd62447: out <= 16'hFF80;
    16'd62448: out <= 16'h01CB;    16'd62449: out <= 16'h0410;    16'd62450: out <= 16'h020B;    16'd62451: out <= 16'h086B;
    16'd62452: out <= 16'h03E7;    16'd62453: out <= 16'hFE3B;    16'd62454: out <= 16'hF5F2;    16'd62455: out <= 16'h0472;
    16'd62456: out <= 16'hFF73;    16'd62457: out <= 16'h02A6;    16'd62458: out <= 16'hFD40;    16'd62459: out <= 16'hFAE0;
    16'd62460: out <= 16'hFD6A;    16'd62461: out <= 16'h0680;    16'd62462: out <= 16'hFF03;    16'd62463: out <= 16'hFBBF;
    16'd62464: out <= 16'h0043;    16'd62465: out <= 16'hFA64;    16'd62466: out <= 16'h04D9;    16'd62467: out <= 16'hFBF0;
    16'd62468: out <= 16'hFF33;    16'd62469: out <= 16'hFDC9;    16'd62470: out <= 16'h04EA;    16'd62471: out <= 16'hF704;
    16'd62472: out <= 16'h0573;    16'd62473: out <= 16'h0171;    16'd62474: out <= 16'hFFCD;    16'd62475: out <= 16'hFA3D;
    16'd62476: out <= 16'hF5A7;    16'd62477: out <= 16'h02C1;    16'd62478: out <= 16'h06BA;    16'd62479: out <= 16'hFF48;
    16'd62480: out <= 16'hFCAA;    16'd62481: out <= 16'hFF5C;    16'd62482: out <= 16'h085A;    16'd62483: out <= 16'hF9E8;
    16'd62484: out <= 16'h044D;    16'd62485: out <= 16'hFF20;    16'd62486: out <= 16'h0323;    16'd62487: out <= 16'h02B7;
    16'd62488: out <= 16'hFF1D;    16'd62489: out <= 16'hFE9D;    16'd62490: out <= 16'h019D;    16'd62491: out <= 16'h03DA;
    16'd62492: out <= 16'hFEF7;    16'd62493: out <= 16'h051E;    16'd62494: out <= 16'h0614;    16'd62495: out <= 16'hFB62;
    16'd62496: out <= 16'hFBC5;    16'd62497: out <= 16'hFFD5;    16'd62498: out <= 16'hFCA0;    16'd62499: out <= 16'hFDB5;
    16'd62500: out <= 16'hF816;    16'd62501: out <= 16'hFA17;    16'd62502: out <= 16'hFA17;    16'd62503: out <= 16'hFD69;
    16'd62504: out <= 16'h0107;    16'd62505: out <= 16'hFE9E;    16'd62506: out <= 16'h0451;    16'd62507: out <= 16'hFAEA;
    16'd62508: out <= 16'h026B;    16'd62509: out <= 16'h00F8;    16'd62510: out <= 16'h006A;    16'd62511: out <= 16'h05D4;
    16'd62512: out <= 16'hFBF6;    16'd62513: out <= 16'h011E;    16'd62514: out <= 16'h01BB;    16'd62515: out <= 16'h01DA;
    16'd62516: out <= 16'h0A4C;    16'd62517: out <= 16'h03B1;    16'd62518: out <= 16'h06D8;    16'd62519: out <= 16'h0720;
    16'd62520: out <= 16'h0500;    16'd62521: out <= 16'h061C;    16'd62522: out <= 16'h0CDD;    16'd62523: out <= 16'h0652;
    16'd62524: out <= 16'h02E1;    16'd62525: out <= 16'h069F;    16'd62526: out <= 16'h082D;    16'd62527: out <= 16'hFFFD;
    16'd62528: out <= 16'h086C;    16'd62529: out <= 16'h01A7;    16'd62530: out <= 16'h019E;    16'd62531: out <= 16'h0D1B;
    16'd62532: out <= 16'h0739;    16'd62533: out <= 16'hFD17;    16'd62534: out <= 16'h01B0;    16'd62535: out <= 16'h0981;
    16'd62536: out <= 16'h038A;    16'd62537: out <= 16'h0471;    16'd62538: out <= 16'h0290;    16'd62539: out <= 16'h0239;
    16'd62540: out <= 16'h0C71;    16'd62541: out <= 16'h03A8;    16'd62542: out <= 16'h08CC;    16'd62543: out <= 16'h0681;
    16'd62544: out <= 16'h0367;    16'd62545: out <= 16'hFF0E;    16'd62546: out <= 16'h063D;    16'd62547: out <= 16'h0079;
    16'd62548: out <= 16'h048A;    16'd62549: out <= 16'hFF41;    16'd62550: out <= 16'h05F8;    16'd62551: out <= 16'hFD91;
    16'd62552: out <= 16'hFD4D;    16'd62553: out <= 16'h020E;    16'd62554: out <= 16'h006A;    16'd62555: out <= 16'hF648;
    16'd62556: out <= 16'h03FB;    16'd62557: out <= 16'hFF73;    16'd62558: out <= 16'hFA96;    16'd62559: out <= 16'h0317;
    16'd62560: out <= 16'h000E;    16'd62561: out <= 16'hFF05;    16'd62562: out <= 16'h005E;    16'd62563: out <= 16'hFCF1;
    16'd62564: out <= 16'hFDA4;    16'd62565: out <= 16'h00B8;    16'd62566: out <= 16'h03D5;    16'd62567: out <= 16'h02B6;
    16'd62568: out <= 16'h0060;    16'd62569: out <= 16'hFB5E;    16'd62570: out <= 16'h0102;    16'd62571: out <= 16'h071D;
    16'd62572: out <= 16'h0189;    16'd62573: out <= 16'h01FD;    16'd62574: out <= 16'h01AD;    16'd62575: out <= 16'hF8F9;
    16'd62576: out <= 16'h00EE;    16'd62577: out <= 16'hFCAB;    16'd62578: out <= 16'hFE63;    16'd62579: out <= 16'h012B;
    16'd62580: out <= 16'h00AA;    16'd62581: out <= 16'hFCF6;    16'd62582: out <= 16'h05B3;    16'd62583: out <= 16'hFC59;
    16'd62584: out <= 16'hFE87;    16'd62585: out <= 16'hFC38;    16'd62586: out <= 16'h03D1;    16'd62587: out <= 16'h0AC9;
    16'd62588: out <= 16'hFBB5;    16'd62589: out <= 16'h0172;    16'd62590: out <= 16'hFC51;    16'd62591: out <= 16'hFB9E;
    16'd62592: out <= 16'hF657;    16'd62593: out <= 16'h067E;    16'd62594: out <= 16'h0159;    16'd62595: out <= 16'hFF08;
    16'd62596: out <= 16'hFE72;    16'd62597: out <= 16'hFBBF;    16'd62598: out <= 16'hF9A1;    16'd62599: out <= 16'hFBA0;
    16'd62600: out <= 16'hFB3B;    16'd62601: out <= 16'h0470;    16'd62602: out <= 16'hFF39;    16'd62603: out <= 16'h05F5;
    16'd62604: out <= 16'hFE27;    16'd62605: out <= 16'hFEBC;    16'd62606: out <= 16'hFAD3;    16'd62607: out <= 16'hFCAA;
    16'd62608: out <= 16'hFF17;    16'd62609: out <= 16'hFF51;    16'd62610: out <= 16'h027A;    16'd62611: out <= 16'hFC9F;
    16'd62612: out <= 16'h0324;    16'd62613: out <= 16'h015A;    16'd62614: out <= 16'hFDCD;    16'd62615: out <= 16'hFED2;
    16'd62616: out <= 16'h054C;    16'd62617: out <= 16'hFF65;    16'd62618: out <= 16'hFA28;    16'd62619: out <= 16'h053F;
    16'd62620: out <= 16'h02B6;    16'd62621: out <= 16'hFC0A;    16'd62622: out <= 16'h0382;    16'd62623: out <= 16'h016B;
    16'd62624: out <= 16'h0195;    16'd62625: out <= 16'hFDC3;    16'd62626: out <= 16'h0122;    16'd62627: out <= 16'h044E;
    16'd62628: out <= 16'h07CA;    16'd62629: out <= 16'hFF95;    16'd62630: out <= 16'h0ACC;    16'd62631: out <= 16'h02D8;
    16'd62632: out <= 16'h07D2;    16'd62633: out <= 16'h0495;    16'd62634: out <= 16'h0818;    16'd62635: out <= 16'h02A0;
    16'd62636: out <= 16'h0558;    16'd62637: out <= 16'h00CD;    16'd62638: out <= 16'h051C;    16'd62639: out <= 16'hFE96;
    16'd62640: out <= 16'h0690;    16'd62641: out <= 16'h0474;    16'd62642: out <= 16'hFF01;    16'd62643: out <= 16'hFCEB;
    16'd62644: out <= 16'h0B99;    16'd62645: out <= 16'h06D2;    16'd62646: out <= 16'h0713;    16'd62647: out <= 16'h085E;
    16'd62648: out <= 16'h02E5;    16'd62649: out <= 16'h0435;    16'd62650: out <= 16'h0D0B;    16'd62651: out <= 16'hFF6E;
    16'd62652: out <= 16'h072B;    16'd62653: out <= 16'h0535;    16'd62654: out <= 16'h008C;    16'd62655: out <= 16'h0325;
    16'd62656: out <= 16'hFEFC;    16'd62657: out <= 16'h0010;    16'd62658: out <= 16'h0461;    16'd62659: out <= 16'h0531;
    16'd62660: out <= 16'hFD8B;    16'd62661: out <= 16'h05A3;    16'd62662: out <= 16'hFDA7;    16'd62663: out <= 16'hFB7A;
    16'd62664: out <= 16'h019A;    16'd62665: out <= 16'hFF2F;    16'd62666: out <= 16'h07C8;    16'd62667: out <= 16'hFCC0;
    16'd62668: out <= 16'h04F0;    16'd62669: out <= 16'h003E;    16'd62670: out <= 16'h02D8;    16'd62671: out <= 16'h0151;
    16'd62672: out <= 16'h04DF;    16'd62673: out <= 16'h057F;    16'd62674: out <= 16'hF980;    16'd62675: out <= 16'hFE27;
    16'd62676: out <= 16'h01A8;    16'd62677: out <= 16'hF751;    16'd62678: out <= 16'h034F;    16'd62679: out <= 16'h0829;
    16'd62680: out <= 16'hFCFB;    16'd62681: out <= 16'h020D;    16'd62682: out <= 16'h035C;    16'd62683: out <= 16'hF37D;
    16'd62684: out <= 16'h012D;    16'd62685: out <= 16'h0200;    16'd62686: out <= 16'h0027;    16'd62687: out <= 16'h01CB;
    16'd62688: out <= 16'hF605;    16'd62689: out <= 16'h05A2;    16'd62690: out <= 16'h0075;    16'd62691: out <= 16'h00D0;
    16'd62692: out <= 16'h0117;    16'd62693: out <= 16'hFCAF;    16'd62694: out <= 16'h03EF;    16'd62695: out <= 16'h0242;
    16'd62696: out <= 16'h046A;    16'd62697: out <= 16'hFB93;    16'd62698: out <= 16'hFF66;    16'd62699: out <= 16'hFE9C;
    16'd62700: out <= 16'h023B;    16'd62701: out <= 16'hFB3F;    16'd62702: out <= 16'h04F6;    16'd62703: out <= 16'h0372;
    16'd62704: out <= 16'hFF4E;    16'd62705: out <= 16'hFFD6;    16'd62706: out <= 16'hFEE7;    16'd62707: out <= 16'hFD6D;
    16'd62708: out <= 16'h0048;    16'd62709: out <= 16'h0279;    16'd62710: out <= 16'h0416;    16'd62711: out <= 16'hFAD4;
    16'd62712: out <= 16'h00C7;    16'd62713: out <= 16'hFF36;    16'd62714: out <= 16'hFC60;    16'd62715: out <= 16'h01DD;
    16'd62716: out <= 16'hFC3E;    16'd62717: out <= 16'h016C;    16'd62718: out <= 16'h010B;    16'd62719: out <= 16'hFC79;
    16'd62720: out <= 16'h04C6;    16'd62721: out <= 16'h03E1;    16'd62722: out <= 16'h076A;    16'd62723: out <= 16'h00BC;
    16'd62724: out <= 16'hFF28;    16'd62725: out <= 16'hFE49;    16'd62726: out <= 16'h0331;    16'd62727: out <= 16'h0361;
    16'd62728: out <= 16'hFC76;    16'd62729: out <= 16'h02FF;    16'd62730: out <= 16'hFB90;    16'd62731: out <= 16'hFE56;
    16'd62732: out <= 16'hFAE1;    16'd62733: out <= 16'hFF6B;    16'd62734: out <= 16'h0901;    16'd62735: out <= 16'h0116;
    16'd62736: out <= 16'h0567;    16'd62737: out <= 16'h0734;    16'd62738: out <= 16'h0435;    16'd62739: out <= 16'h0429;
    16'd62740: out <= 16'h00E0;    16'd62741: out <= 16'h00C2;    16'd62742: out <= 16'hFCBB;    16'd62743: out <= 16'hFEC7;
    16'd62744: out <= 16'hFEC1;    16'd62745: out <= 16'hF7DD;    16'd62746: out <= 16'h009E;    16'd62747: out <= 16'h0794;
    16'd62748: out <= 16'h0398;    16'd62749: out <= 16'hFFA9;    16'd62750: out <= 16'h0289;    16'd62751: out <= 16'h06C8;
    16'd62752: out <= 16'hFF23;    16'd62753: out <= 16'h01EF;    16'd62754: out <= 16'h02B9;    16'd62755: out <= 16'h0217;
    16'd62756: out <= 16'h04CB;    16'd62757: out <= 16'h027C;    16'd62758: out <= 16'hFC68;    16'd62759: out <= 16'h05C6;
    16'd62760: out <= 16'hFE31;    16'd62761: out <= 16'hFB32;    16'd62762: out <= 16'h07FA;    16'd62763: out <= 16'h0068;
    16'd62764: out <= 16'h04CD;    16'd62765: out <= 16'h0BC6;    16'd62766: out <= 16'h01BB;    16'd62767: out <= 16'h0935;
    16'd62768: out <= 16'h0118;    16'd62769: out <= 16'h01CC;    16'd62770: out <= 16'h0603;    16'd62771: out <= 16'h04F8;
    16'd62772: out <= 16'h0308;    16'd62773: out <= 16'h046A;    16'd62774: out <= 16'h062D;    16'd62775: out <= 16'h05D0;
    16'd62776: out <= 16'h0120;    16'd62777: out <= 16'hFD25;    16'd62778: out <= 16'h0804;    16'd62779: out <= 16'h04E6;
    16'd62780: out <= 16'h0698;    16'd62781: out <= 16'hFD2C;    16'd62782: out <= 16'h0655;    16'd62783: out <= 16'h0675;
    16'd62784: out <= 16'hFF3D;    16'd62785: out <= 16'h0A24;    16'd62786: out <= 16'h0420;    16'd62787: out <= 16'h0D2A;
    16'd62788: out <= 16'h0840;    16'd62789: out <= 16'h01DF;    16'd62790: out <= 16'hFF84;    16'd62791: out <= 16'h0B10;
    16'd62792: out <= 16'hFD05;    16'd62793: out <= 16'h0219;    16'd62794: out <= 16'h0145;    16'd62795: out <= 16'h0274;
    16'd62796: out <= 16'h00BA;    16'd62797: out <= 16'h0077;    16'd62798: out <= 16'hFF55;    16'd62799: out <= 16'h0991;
    16'd62800: out <= 16'h066D;    16'd62801: out <= 16'hFFE6;    16'd62802: out <= 16'h01FF;    16'd62803: out <= 16'h008C;
    16'd62804: out <= 16'h03B3;    16'd62805: out <= 16'hFEE6;    16'd62806: out <= 16'hFB5D;    16'd62807: out <= 16'h0472;
    16'd62808: out <= 16'h02CC;    16'd62809: out <= 16'hFD80;    16'd62810: out <= 16'h02A6;    16'd62811: out <= 16'h0176;
    16'd62812: out <= 16'h00FD;    16'd62813: out <= 16'hFE94;    16'd62814: out <= 16'hFD18;    16'd62815: out <= 16'h0267;
    16'd62816: out <= 16'h0076;    16'd62817: out <= 16'hFD14;    16'd62818: out <= 16'h0227;    16'd62819: out <= 16'hFC5C;
    16'd62820: out <= 16'hFE9A;    16'd62821: out <= 16'hFF1C;    16'd62822: out <= 16'h0156;    16'd62823: out <= 16'hFFC8;
    16'd62824: out <= 16'hFCA5;    16'd62825: out <= 16'h078F;    16'd62826: out <= 16'h064E;    16'd62827: out <= 16'h041C;
    16'd62828: out <= 16'hFCF3;    16'd62829: out <= 16'hFD4D;    16'd62830: out <= 16'hFDB5;    16'd62831: out <= 16'h009D;
    16'd62832: out <= 16'h0231;    16'd62833: out <= 16'hFAA0;    16'd62834: out <= 16'hFF01;    16'd62835: out <= 16'hFEC0;
    16'd62836: out <= 16'hFCDF;    16'd62837: out <= 16'hFF24;    16'd62838: out <= 16'hFEBA;    16'd62839: out <= 16'hFF8F;
    16'd62840: out <= 16'hFD44;    16'd62841: out <= 16'hFF64;    16'd62842: out <= 16'hFE9E;    16'd62843: out <= 16'h00C2;
    16'd62844: out <= 16'hFFAC;    16'd62845: out <= 16'hFAEA;    16'd62846: out <= 16'h0BD5;    16'd62847: out <= 16'h0488;
    16'd62848: out <= 16'h004E;    16'd62849: out <= 16'hF8A3;    16'd62850: out <= 16'hFFD4;    16'd62851: out <= 16'h0364;
    16'd62852: out <= 16'h020F;    16'd62853: out <= 16'hFDA9;    16'd62854: out <= 16'hFE82;    16'd62855: out <= 16'hFB78;
    16'd62856: out <= 16'hFFC5;    16'd62857: out <= 16'h000E;    16'd62858: out <= 16'hFE3D;    16'd62859: out <= 16'hFABD;
    16'd62860: out <= 16'h0738;    16'd62861: out <= 16'hFE6E;    16'd62862: out <= 16'hFE37;    16'd62863: out <= 16'h001B;
    16'd62864: out <= 16'h00FA;    16'd62865: out <= 16'hFDA2;    16'd62866: out <= 16'h023A;    16'd62867: out <= 16'h00D6;
    16'd62868: out <= 16'h04FC;    16'd62869: out <= 16'hFE4B;    16'd62870: out <= 16'hF681;    16'd62871: out <= 16'hFB09;
    16'd62872: out <= 16'hFED9;    16'd62873: out <= 16'h01E7;    16'd62874: out <= 16'hFA91;    16'd62875: out <= 16'h03CA;
    16'd62876: out <= 16'hFD6F;    16'd62877: out <= 16'h022E;    16'd62878: out <= 16'h09A5;    16'd62879: out <= 16'h000B;
    16'd62880: out <= 16'h05B5;    16'd62881: out <= 16'hF858;    16'd62882: out <= 16'h0550;    16'd62883: out <= 16'hFD1B;
    16'd62884: out <= 16'hFD98;    16'd62885: out <= 16'h0BD4;    16'd62886: out <= 16'h0858;    16'd62887: out <= 16'h06FC;
    16'd62888: out <= 16'h0313;    16'd62889: out <= 16'h054A;    16'd62890: out <= 16'h051E;    16'd62891: out <= 16'h00C3;
    16'd62892: out <= 16'hFD0A;    16'd62893: out <= 16'h0263;    16'd62894: out <= 16'hFDEA;    16'd62895: out <= 16'h03B4;
    16'd62896: out <= 16'hFE7B;    16'd62897: out <= 16'h08EC;    16'd62898: out <= 16'h00C5;    16'd62899: out <= 16'h0464;
    16'd62900: out <= 16'h0320;    16'd62901: out <= 16'hFF9D;    16'd62902: out <= 16'h011F;    16'd62903: out <= 16'h062F;
    16'd62904: out <= 16'h0194;    16'd62905: out <= 16'hFCE1;    16'd62906: out <= 16'h044E;    16'd62907: out <= 16'hFE9B;
    16'd62908: out <= 16'hFD9F;    16'd62909: out <= 16'h00D2;    16'd62910: out <= 16'h0267;    16'd62911: out <= 16'h08B0;
    16'd62912: out <= 16'h03FB;    16'd62913: out <= 16'h0486;    16'd62914: out <= 16'h00FD;    16'd62915: out <= 16'h06B6;
    16'd62916: out <= 16'h007D;    16'd62917: out <= 16'h0408;    16'd62918: out <= 16'h061F;    16'd62919: out <= 16'h0323;
    16'd62920: out <= 16'h027F;    16'd62921: out <= 16'h053F;    16'd62922: out <= 16'h0082;    16'd62923: out <= 16'h03A4;
    16'd62924: out <= 16'h02D3;    16'd62925: out <= 16'hFAC1;    16'd62926: out <= 16'h0303;    16'd62927: out <= 16'hFAD2;
    16'd62928: out <= 16'h072C;    16'd62929: out <= 16'h03C5;    16'd62930: out <= 16'hFF30;    16'd62931: out <= 16'hFAE0;
    16'd62932: out <= 16'hF6CE;    16'd62933: out <= 16'h039E;    16'd62934: out <= 16'h00CA;    16'd62935: out <= 16'h0399;
    16'd62936: out <= 16'hFD5E;    16'd62937: out <= 16'hFBAF;    16'd62938: out <= 16'hFFC9;    16'd62939: out <= 16'hFF51;
    16'd62940: out <= 16'hF8C9;    16'd62941: out <= 16'h0275;    16'd62942: out <= 16'h0312;    16'd62943: out <= 16'hFDFE;
    16'd62944: out <= 16'hFC1F;    16'd62945: out <= 16'hFF53;    16'd62946: out <= 16'hFFC1;    16'd62947: out <= 16'h00ED;
    16'd62948: out <= 16'h0680;    16'd62949: out <= 16'h085F;    16'd62950: out <= 16'h02FB;    16'd62951: out <= 16'hFD8F;
    16'd62952: out <= 16'h03E8;    16'd62953: out <= 16'h08F7;    16'd62954: out <= 16'hFCC3;    16'd62955: out <= 16'h02AC;
    16'd62956: out <= 16'h060D;    16'd62957: out <= 16'h038A;    16'd62958: out <= 16'hFA72;    16'd62959: out <= 16'h0491;
    16'd62960: out <= 16'hFF96;    16'd62961: out <= 16'hFF3B;    16'd62962: out <= 16'hFDC3;    16'd62963: out <= 16'hFDAA;
    16'd62964: out <= 16'h0255;    16'd62965: out <= 16'h042E;    16'd62966: out <= 16'h0000;    16'd62967: out <= 16'h0004;
    16'd62968: out <= 16'hFEFC;    16'd62969: out <= 16'h00EE;    16'd62970: out <= 16'hFB07;    16'd62971: out <= 16'hFE9B;
    16'd62972: out <= 16'hFEEB;    16'd62973: out <= 16'hF7D3;    16'd62974: out <= 16'hF949;    16'd62975: out <= 16'h017C;
    16'd62976: out <= 16'hFB4C;    16'd62977: out <= 16'h015B;    16'd62978: out <= 16'hFE90;    16'd62979: out <= 16'h03FA;
    16'd62980: out <= 16'hFBBE;    16'd62981: out <= 16'h0994;    16'd62982: out <= 16'h0240;    16'd62983: out <= 16'hFDF4;
    16'd62984: out <= 16'hFEA4;    16'd62985: out <= 16'h062F;    16'd62986: out <= 16'h0A2C;    16'd62987: out <= 16'hFCFE;
    16'd62988: out <= 16'h03FB;    16'd62989: out <= 16'hFC3C;    16'd62990: out <= 16'hFE2A;    16'd62991: out <= 16'hFF37;
    16'd62992: out <= 16'h049E;    16'd62993: out <= 16'hFF6D;    16'd62994: out <= 16'h02D1;    16'd62995: out <= 16'h01AF;
    16'd62996: out <= 16'hFFFA;    16'd62997: out <= 16'hFDD5;    16'd62998: out <= 16'hFDC2;    16'd62999: out <= 16'h0D02;
    16'd63000: out <= 16'h027F;    16'd63001: out <= 16'h03B5;    16'd63002: out <= 16'h001C;    16'd63003: out <= 16'h0596;
    16'd63004: out <= 16'h095B;    16'd63005: out <= 16'h0146;    16'd63006: out <= 16'hF9F3;    16'd63007: out <= 16'h04BB;
    16'd63008: out <= 16'hFB8D;    16'd63009: out <= 16'hFE8F;    16'd63010: out <= 16'h04E0;    16'd63011: out <= 16'hFF27;
    16'd63012: out <= 16'h0537;    16'd63013: out <= 16'h0074;    16'd63014: out <= 16'h0284;    16'd63015: out <= 16'h00F1;
    16'd63016: out <= 16'h03B1;    16'd63017: out <= 16'h007C;    16'd63018: out <= 16'hFF95;    16'd63019: out <= 16'h0D4F;
    16'd63020: out <= 16'h0298;    16'd63021: out <= 16'h030B;    16'd63022: out <= 16'h0659;    16'd63023: out <= 16'h040E;
    16'd63024: out <= 16'hFE99;    16'd63025: out <= 16'h04F5;    16'd63026: out <= 16'h02CF;    16'd63027: out <= 16'h034C;
    16'd63028: out <= 16'h091E;    16'd63029: out <= 16'h07E3;    16'd63030: out <= 16'h0547;    16'd63031: out <= 16'h05F2;
    16'd63032: out <= 16'h0579;    16'd63033: out <= 16'hFDBE;    16'd63034: out <= 16'h009F;    16'd63035: out <= 16'hFF1B;
    16'd63036: out <= 16'h058F;    16'd63037: out <= 16'h02C6;    16'd63038: out <= 16'h01CB;    16'd63039: out <= 16'h0AD6;
    16'd63040: out <= 16'hFDFD;    16'd63041: out <= 16'h05D1;    16'd63042: out <= 16'h03BF;    16'd63043: out <= 16'h0429;
    16'd63044: out <= 16'h075B;    16'd63045: out <= 16'h00AD;    16'd63046: out <= 16'h0721;    16'd63047: out <= 16'h05C1;
    16'd63048: out <= 16'h013A;    16'd63049: out <= 16'h0663;    16'd63050: out <= 16'h0365;    16'd63051: out <= 16'h0AC1;
    16'd63052: out <= 16'h078D;    16'd63053: out <= 16'h054F;    16'd63054: out <= 16'h0215;    16'd63055: out <= 16'h0799;
    16'd63056: out <= 16'h05D6;    16'd63057: out <= 16'h03E6;    16'd63058: out <= 16'h0431;    16'd63059: out <= 16'h0811;
    16'd63060: out <= 16'h049C;    16'd63061: out <= 16'h0627;    16'd63062: out <= 16'hFF60;    16'd63063: out <= 16'h0028;
    16'd63064: out <= 16'hFD3F;    16'd63065: out <= 16'h000D;    16'd63066: out <= 16'h0572;    16'd63067: out <= 16'hFF6A;
    16'd63068: out <= 16'hFE10;    16'd63069: out <= 16'hFB72;    16'd63070: out <= 16'h00E8;    16'd63071: out <= 16'hFE39;
    16'd63072: out <= 16'h0208;    16'd63073: out <= 16'h0101;    16'd63074: out <= 16'h04E8;    16'd63075: out <= 16'hFC6E;
    16'd63076: out <= 16'hFC4F;    16'd63077: out <= 16'hFED1;    16'd63078: out <= 16'h06AE;    16'd63079: out <= 16'h0217;
    16'd63080: out <= 16'hFA33;    16'd63081: out <= 16'h0062;    16'd63082: out <= 16'hFE4C;    16'd63083: out <= 16'h03C7;
    16'd63084: out <= 16'hFF1B;    16'd63085: out <= 16'h0025;    16'd63086: out <= 16'hFFBE;    16'd63087: out <= 16'hFD17;
    16'd63088: out <= 16'h0398;    16'd63089: out <= 16'hFF35;    16'd63090: out <= 16'hFDE2;    16'd63091: out <= 16'hFEDA;
    16'd63092: out <= 16'hFAEF;    16'd63093: out <= 16'hFAB5;    16'd63094: out <= 16'h0903;    16'd63095: out <= 16'h0221;
    16'd63096: out <= 16'hF96D;    16'd63097: out <= 16'hFE1B;    16'd63098: out <= 16'h023A;    16'd63099: out <= 16'hFD52;
    16'd63100: out <= 16'hF987;    16'd63101: out <= 16'hFD39;    16'd63102: out <= 16'h01C9;    16'd63103: out <= 16'h0142;
    16'd63104: out <= 16'hFFA8;    16'd63105: out <= 16'hFCD1;    16'd63106: out <= 16'h028D;    16'd63107: out <= 16'h0549;
    16'd63108: out <= 16'hFF33;    16'd63109: out <= 16'hF9F7;    16'd63110: out <= 16'hFCA3;    16'd63111: out <= 16'hFC8F;
    16'd63112: out <= 16'h00B4;    16'd63113: out <= 16'hF794;    16'd63114: out <= 16'h02BB;    16'd63115: out <= 16'h0342;
    16'd63116: out <= 16'hFC5E;    16'd63117: out <= 16'h0673;    16'd63118: out <= 16'h09AB;    16'd63119: out <= 16'hFEF5;
    16'd63120: out <= 16'hFB12;    16'd63121: out <= 16'hF914;    16'd63122: out <= 16'h00F9;    16'd63123: out <= 16'hFC20;
    16'd63124: out <= 16'hFEBC;    16'd63125: out <= 16'h0004;    16'd63126: out <= 16'hFD1B;    16'd63127: out <= 16'hFCB4;
    16'd63128: out <= 16'hFB4B;    16'd63129: out <= 16'h06E4;    16'd63130: out <= 16'hFA6C;    16'd63131: out <= 16'h02A6;
    16'd63132: out <= 16'hFEC8;    16'd63133: out <= 16'h012C;    16'd63134: out <= 16'h00D8;    16'd63135: out <= 16'h0140;
    16'd63136: out <= 16'hFDB4;    16'd63137: out <= 16'hFD37;    16'd63138: out <= 16'h03CB;    16'd63139: out <= 16'h025E;
    16'd63140: out <= 16'h01CA;    16'd63141: out <= 16'h06E6;    16'd63142: out <= 16'h0491;    16'd63143: out <= 16'h0566;
    16'd63144: out <= 16'h0642;    16'd63145: out <= 16'h0088;    16'd63146: out <= 16'h01DB;    16'd63147: out <= 16'hFF0E;
    16'd63148: out <= 16'h0007;    16'd63149: out <= 16'hF8FC;    16'd63150: out <= 16'h070A;    16'd63151: out <= 16'h03EC;
    16'd63152: out <= 16'h0185;    16'd63153: out <= 16'h01FB;    16'd63154: out <= 16'h0BBF;    16'd63155: out <= 16'h035C;
    16'd63156: out <= 16'h0CB1;    16'd63157: out <= 16'h07DC;    16'd63158: out <= 16'h0348;    16'd63159: out <= 16'h0448;
    16'd63160: out <= 16'h0356;    16'd63161: out <= 16'hFDCA;    16'd63162: out <= 16'h0B06;    16'd63163: out <= 16'hFC3E;
    16'd63164: out <= 16'h08DC;    16'd63165: out <= 16'h09EB;    16'd63166: out <= 16'h03FD;    16'd63167: out <= 16'h0DFF;
    16'd63168: out <= 16'h05D5;    16'd63169: out <= 16'hFF92;    16'd63170: out <= 16'h065D;    16'd63171: out <= 16'h00E8;
    16'd63172: out <= 16'h0049;    16'd63173: out <= 16'h08B3;    16'd63174: out <= 16'hFD01;    16'd63175: out <= 16'hF687;
    16'd63176: out <= 16'hF513;    16'd63177: out <= 16'h015E;    16'd63178: out <= 16'hFD7A;    16'd63179: out <= 16'hFD3A;
    16'd63180: out <= 16'hFBC0;    16'd63181: out <= 16'hF976;    16'd63182: out <= 16'h018D;    16'd63183: out <= 16'h054A;
    16'd63184: out <= 16'hFBF0;    16'd63185: out <= 16'h0316;    16'd63186: out <= 16'hFE6A;    16'd63187: out <= 16'h0615;
    16'd63188: out <= 16'h0021;    16'd63189: out <= 16'hFC62;    16'd63190: out <= 16'hFF7D;    16'd63191: out <= 16'h0525;
    16'd63192: out <= 16'h02D8;    16'd63193: out <= 16'hFD1F;    16'd63194: out <= 16'hF855;    16'd63195: out <= 16'hFE2F;
    16'd63196: out <= 16'hFF0F;    16'd63197: out <= 16'h013B;    16'd63198: out <= 16'h0447;    16'd63199: out <= 16'h01B7;
    16'd63200: out <= 16'hFF7D;    16'd63201: out <= 16'hFFBB;    16'd63202: out <= 16'h0303;    16'd63203: out <= 16'h0382;
    16'd63204: out <= 16'hFC32;    16'd63205: out <= 16'hFF13;    16'd63206: out <= 16'h05D6;    16'd63207: out <= 16'hFF24;
    16'd63208: out <= 16'h0166;    16'd63209: out <= 16'h0443;    16'd63210: out <= 16'hF64F;    16'd63211: out <= 16'h0734;
    16'd63212: out <= 16'h02B9;    16'd63213: out <= 16'h008D;    16'd63214: out <= 16'hFE8D;    16'd63215: out <= 16'hFE34;
    16'd63216: out <= 16'hFEE5;    16'd63217: out <= 16'hFEFE;    16'd63218: out <= 16'hF4D0;    16'd63219: out <= 16'h05B9;
    16'd63220: out <= 16'hFF79;    16'd63221: out <= 16'hFCB9;    16'd63222: out <= 16'h0ACE;    16'd63223: out <= 16'h00BF;
    16'd63224: out <= 16'hFAF6;    16'd63225: out <= 16'h0111;    16'd63226: out <= 16'h03D4;    16'd63227: out <= 16'h0550;
    16'd63228: out <= 16'hFB57;    16'd63229: out <= 16'hFF4A;    16'd63230: out <= 16'h0264;    16'd63231: out <= 16'hFF70;
    16'd63232: out <= 16'h067B;    16'd63233: out <= 16'hFF96;    16'd63234: out <= 16'hFDC4;    16'd63235: out <= 16'hFFC7;
    16'd63236: out <= 16'h05F6;    16'd63237: out <= 16'h00B6;    16'd63238: out <= 16'hFDD9;    16'd63239: out <= 16'hFC73;
    16'd63240: out <= 16'h0558;    16'd63241: out <= 16'hFDD8;    16'd63242: out <= 16'hFDC0;    16'd63243: out <= 16'h053D;
    16'd63244: out <= 16'h04CC;    16'd63245: out <= 16'hFEF0;    16'd63246: out <= 16'hFFDF;    16'd63247: out <= 16'hFDA2;
    16'd63248: out <= 16'hFF10;    16'd63249: out <= 16'hFF95;    16'd63250: out <= 16'h0502;    16'd63251: out <= 16'hFBE8;
    16'd63252: out <= 16'h02C5;    16'd63253: out <= 16'hFD43;    16'd63254: out <= 16'hFC83;    16'd63255: out <= 16'hFC1D;
    16'd63256: out <= 16'h06CD;    16'd63257: out <= 16'hFDB8;    16'd63258: out <= 16'hFD36;    16'd63259: out <= 16'hF94C;
    16'd63260: out <= 16'hF93C;    16'd63261: out <= 16'h0294;    16'd63262: out <= 16'h0307;    16'd63263: out <= 16'hF903;
    16'd63264: out <= 16'h0016;    16'd63265: out <= 16'hFCA0;    16'd63266: out <= 16'h0D41;    16'd63267: out <= 16'h04AC;
    16'd63268: out <= 16'h0BD7;    16'd63269: out <= 16'hFD55;    16'd63270: out <= 16'h0178;    16'd63271: out <= 16'hFA7A;
    16'd63272: out <= 16'h01C8;    16'd63273: out <= 16'hFBA0;    16'd63274: out <= 16'h0679;    16'd63275: out <= 16'hFCD7;
    16'd63276: out <= 16'h00DF;    16'd63277: out <= 16'h03FF;    16'd63278: out <= 16'h06E6;    16'd63279: out <= 16'hFF11;
    16'd63280: out <= 16'h022D;    16'd63281: out <= 16'h0AA4;    16'd63282: out <= 16'h0523;    16'd63283: out <= 16'h0A61;
    16'd63284: out <= 16'h04F3;    16'd63285: out <= 16'h0823;    16'd63286: out <= 16'h045D;    16'd63287: out <= 16'h039A;
    16'd63288: out <= 16'h0927;    16'd63289: out <= 16'h0421;    16'd63290: out <= 16'hFE67;    16'd63291: out <= 16'h025E;
    16'd63292: out <= 16'hF948;    16'd63293: out <= 16'h0AD6;    16'd63294: out <= 16'h02E8;    16'd63295: out <= 16'h0819;
    16'd63296: out <= 16'h0863;    16'd63297: out <= 16'h0522;    16'd63298: out <= 16'h011A;    16'd63299: out <= 16'h02D3;
    16'd63300: out <= 16'hFF9E;    16'd63301: out <= 16'hFE4D;    16'd63302: out <= 16'h07C8;    16'd63303: out <= 16'h07F5;
    16'd63304: out <= 16'hFED5;    16'd63305: out <= 16'h03E1;    16'd63306: out <= 16'h054A;    16'd63307: out <= 16'h0101;
    16'd63308: out <= 16'h035E;    16'd63309: out <= 16'h041E;    16'd63310: out <= 16'h0045;    16'd63311: out <= 16'h079E;
    16'd63312: out <= 16'h0400;    16'd63313: out <= 16'h04C7;    16'd63314: out <= 16'h07E0;    16'd63315: out <= 16'h0049;
    16'd63316: out <= 16'h02A5;    16'd63317: out <= 16'hFEFC;    16'd63318: out <= 16'h09FE;    16'd63319: out <= 16'h0111;
    16'd63320: out <= 16'hF8A3;    16'd63321: out <= 16'h006D;    16'd63322: out <= 16'h0240;    16'd63323: out <= 16'h0194;
    16'd63324: out <= 16'h00E2;    16'd63325: out <= 16'h02BC;    16'd63326: out <= 16'hFB91;    16'd63327: out <= 16'h09B2;
    16'd63328: out <= 16'hFB62;    16'd63329: out <= 16'hFF3B;    16'd63330: out <= 16'h04CE;    16'd63331: out <= 16'hF994;
    16'd63332: out <= 16'hFD11;    16'd63333: out <= 16'hFDEA;    16'd63334: out <= 16'h0AC4;    16'd63335: out <= 16'hFD6E;
    16'd63336: out <= 16'h00C3;    16'd63337: out <= 16'h007F;    16'd63338: out <= 16'h0676;    16'd63339: out <= 16'hFE17;
    16'd63340: out <= 16'hFEF4;    16'd63341: out <= 16'hFFCC;    16'd63342: out <= 16'h0104;    16'd63343: out <= 16'hFB60;
    16'd63344: out <= 16'hFF0D;    16'd63345: out <= 16'hFF7C;    16'd63346: out <= 16'h0239;    16'd63347: out <= 16'h0396;
    16'd63348: out <= 16'h0142;    16'd63349: out <= 16'h03B8;    16'd63350: out <= 16'h02E7;    16'd63351: out <= 16'h02BB;
    16'd63352: out <= 16'h034C;    16'd63353: out <= 16'h005F;    16'd63354: out <= 16'hFD20;    16'd63355: out <= 16'hFD2A;
    16'd63356: out <= 16'hFF9F;    16'd63357: out <= 16'hFE37;    16'd63358: out <= 16'h06C0;    16'd63359: out <= 16'hFC53;
    16'd63360: out <= 16'h03E0;    16'd63361: out <= 16'h0150;    16'd63362: out <= 16'h030D;    16'd63363: out <= 16'hFB5C;
    16'd63364: out <= 16'h0219;    16'd63365: out <= 16'hFECC;    16'd63366: out <= 16'hFE56;    16'd63367: out <= 16'hF557;
    16'd63368: out <= 16'h0174;    16'd63369: out <= 16'h000A;    16'd63370: out <= 16'h0117;    16'd63371: out <= 16'hFC09;
    16'd63372: out <= 16'hFE73;    16'd63373: out <= 16'h0099;    16'd63374: out <= 16'h031C;    16'd63375: out <= 16'hFDFA;
    16'd63376: out <= 16'hFEF2;    16'd63377: out <= 16'hFDB5;    16'd63378: out <= 16'h0012;    16'd63379: out <= 16'h0281;
    16'd63380: out <= 16'h053D;    16'd63381: out <= 16'hFD09;    16'd63382: out <= 16'h05D2;    16'd63383: out <= 16'hFCB4;
    16'd63384: out <= 16'h00D4;    16'd63385: out <= 16'h019E;    16'd63386: out <= 16'hFB32;    16'd63387: out <= 16'hFE45;
    16'd63388: out <= 16'h020E;    16'd63389: out <= 16'h00CE;    16'd63390: out <= 16'h0437;    16'd63391: out <= 16'hFC98;
    16'd63392: out <= 16'h03F2;    16'd63393: out <= 16'h03B4;    16'd63394: out <= 16'h01C0;    16'd63395: out <= 16'h03F2;
    16'd63396: out <= 16'h038B;    16'd63397: out <= 16'h005D;    16'd63398: out <= 16'h02C1;    16'd63399: out <= 16'h0A8B;
    16'd63400: out <= 16'h035E;    16'd63401: out <= 16'h05C7;    16'd63402: out <= 16'h011C;    16'd63403: out <= 16'h05A3;
    16'd63404: out <= 16'hFF44;    16'd63405: out <= 16'h02C0;    16'd63406: out <= 16'h03B5;    16'd63407: out <= 16'h0203;
    16'd63408: out <= 16'h076E;    16'd63409: out <= 16'hFF10;    16'd63410: out <= 16'h06E1;    16'd63411: out <= 16'h0822;
    16'd63412: out <= 16'h0440;    16'd63413: out <= 16'h0231;    16'd63414: out <= 16'h0095;    16'd63415: out <= 16'h01D5;
    16'd63416: out <= 16'hFFC1;    16'd63417: out <= 16'h0226;    16'd63418: out <= 16'h037F;    16'd63419: out <= 16'hFEA5;
    16'd63420: out <= 16'h054C;    16'd63421: out <= 16'h022D;    16'd63422: out <= 16'h0591;    16'd63423: out <= 16'hFE41;
    16'd63424: out <= 16'h028F;    16'd63425: out <= 16'h022A;    16'd63426: out <= 16'h05E6;    16'd63427: out <= 16'h013A;
    16'd63428: out <= 16'h04FF;    16'd63429: out <= 16'h030F;    16'd63430: out <= 16'hFF61;    16'd63431: out <= 16'hFC56;
    16'd63432: out <= 16'h0709;    16'd63433: out <= 16'hFDCF;    16'd63434: out <= 16'hFF59;    16'd63435: out <= 16'h0078;
    16'd63436: out <= 16'hF9C6;    16'd63437: out <= 16'hFBAC;    16'd63438: out <= 16'hF857;    16'd63439: out <= 16'hFC57;
    16'd63440: out <= 16'h036E;    16'd63441: out <= 16'h03E5;    16'd63442: out <= 16'h0492;    16'd63443: out <= 16'h02C8;
    16'd63444: out <= 16'h02BC;    16'd63445: out <= 16'h00BE;    16'd63446: out <= 16'hFE2B;    16'd63447: out <= 16'h06C0;
    16'd63448: out <= 16'h00BD;    16'd63449: out <= 16'hFC46;    16'd63450: out <= 16'hFCD2;    16'd63451: out <= 16'h097B;
    16'd63452: out <= 16'h0361;    16'd63453: out <= 16'hFD3D;    16'd63454: out <= 16'hFCEE;    16'd63455: out <= 16'hFA33;
    16'd63456: out <= 16'h022E;    16'd63457: out <= 16'h017C;    16'd63458: out <= 16'h029A;    16'd63459: out <= 16'h073C;
    16'd63460: out <= 16'h0405;    16'd63461: out <= 16'h02AB;    16'd63462: out <= 16'hF988;    16'd63463: out <= 16'h074A;
    16'd63464: out <= 16'h052B;    16'd63465: out <= 16'h023D;    16'd63466: out <= 16'h008D;    16'd63467: out <= 16'h01FD;
    16'd63468: out <= 16'h0771;    16'd63469: out <= 16'hFD93;    16'd63470: out <= 16'h04E5;    16'd63471: out <= 16'h0440;
    16'd63472: out <= 16'hFF9C;    16'd63473: out <= 16'h02FF;    16'd63474: out <= 16'h0734;    16'd63475: out <= 16'h0194;
    16'd63476: out <= 16'h0260;    16'd63477: out <= 16'h03D0;    16'd63478: out <= 16'h030A;    16'd63479: out <= 16'hFC8A;
    16'd63480: out <= 16'hF680;    16'd63481: out <= 16'h0011;    16'd63482: out <= 16'h00BE;    16'd63483: out <= 16'hFEE5;
    16'd63484: out <= 16'hFAB3;    16'd63485: out <= 16'hFE4D;    16'd63486: out <= 16'h01D5;    16'd63487: out <= 16'h0030;
    16'd63488: out <= 16'h01EB;    16'd63489: out <= 16'hFDDC;    16'd63490: out <= 16'h0186;    16'd63491: out <= 16'h04C1;
    16'd63492: out <= 16'hF67A;    16'd63493: out <= 16'hFBC6;    16'd63494: out <= 16'h0433;    16'd63495: out <= 16'hFAC9;
    16'd63496: out <= 16'hFEBD;    16'd63497: out <= 16'hFEDB;    16'd63498: out <= 16'hFF1F;    16'd63499: out <= 16'h018F;
    16'd63500: out <= 16'hF665;    16'd63501: out <= 16'hFC64;    16'd63502: out <= 16'hFCB2;    16'd63503: out <= 16'h0648;
    16'd63504: out <= 16'h01CC;    16'd63505: out <= 16'hFE13;    16'd63506: out <= 16'h017E;    16'd63507: out <= 16'hFF95;
    16'd63508: out <= 16'hF91B;    16'd63509: out <= 16'hFBC0;    16'd63510: out <= 16'h0300;    16'd63511: out <= 16'hFE49;
    16'd63512: out <= 16'hFE4C;    16'd63513: out <= 16'hFD22;    16'd63514: out <= 16'h01B3;    16'd63515: out <= 16'hFCE6;
    16'd63516: out <= 16'hFEE6;    16'd63517: out <= 16'h00EE;    16'd63518: out <= 16'h01EB;    16'd63519: out <= 16'h06BA;
    16'd63520: out <= 16'h005B;    16'd63521: out <= 16'h006C;    16'd63522: out <= 16'hFC8C;    16'd63523: out <= 16'h00E7;
    16'd63524: out <= 16'h007F;    16'd63525: out <= 16'h0697;    16'd63526: out <= 16'hFE3C;    16'd63527: out <= 16'hF85F;
    16'd63528: out <= 16'hFACE;    16'd63529: out <= 16'hF9CA;    16'd63530: out <= 16'h0195;    16'd63531: out <= 16'h094A;
    16'd63532: out <= 16'h0902;    16'd63533: out <= 16'h0900;    16'd63534: out <= 16'hFDBB;    16'd63535: out <= 16'h0072;
    16'd63536: out <= 16'h04CB;    16'd63537: out <= 16'h024E;    16'd63538: out <= 16'h10FC;    16'd63539: out <= 16'h0A07;
    16'd63540: out <= 16'h00DA;    16'd63541: out <= 16'h011A;    16'd63542: out <= 16'h0447;    16'd63543: out <= 16'h0399;
    16'd63544: out <= 16'h03E8;    16'd63545: out <= 16'h003D;    16'd63546: out <= 16'hFFF2;    16'd63547: out <= 16'h0595;
    16'd63548: out <= 16'h03A3;    16'd63549: out <= 16'h0604;    16'd63550: out <= 16'h03B6;    16'd63551: out <= 16'h01B3;
    16'd63552: out <= 16'h01F2;    16'd63553: out <= 16'h069A;    16'd63554: out <= 16'h035E;    16'd63555: out <= 16'h00F6;
    16'd63556: out <= 16'h0673;    16'd63557: out <= 16'h09C3;    16'd63558: out <= 16'h0383;    16'd63559: out <= 16'h04BE;
    16'd63560: out <= 16'h0BE9;    16'd63561: out <= 16'hFE3E;    16'd63562: out <= 16'h0B77;    16'd63563: out <= 16'h02DB;
    16'd63564: out <= 16'h06B9;    16'd63565: out <= 16'h05FA;    16'd63566: out <= 16'hFD9A;    16'd63567: out <= 16'h02C4;
    16'd63568: out <= 16'h04C6;    16'd63569: out <= 16'h092E;    16'd63570: out <= 16'h0338;    16'd63571: out <= 16'h02EA;
    16'd63572: out <= 16'h03C1;    16'd63573: out <= 16'hFD38;    16'd63574: out <= 16'h0A0C;    16'd63575: out <= 16'hFE85;
    16'd63576: out <= 16'hFE09;    16'd63577: out <= 16'hFFD6;    16'd63578: out <= 16'hF940;    16'd63579: out <= 16'hFEF2;
    16'd63580: out <= 16'hFDB0;    16'd63581: out <= 16'h056F;    16'd63582: out <= 16'h0044;    16'd63583: out <= 16'h0385;
    16'd63584: out <= 16'hFFEE;    16'd63585: out <= 16'hFDC9;    16'd63586: out <= 16'h0226;    16'd63587: out <= 16'hFBD1;
    16'd63588: out <= 16'hFF5B;    16'd63589: out <= 16'h095F;    16'd63590: out <= 16'h07C9;    16'd63591: out <= 16'h042E;
    16'd63592: out <= 16'h04B7;    16'd63593: out <= 16'h0254;    16'd63594: out <= 16'hFD96;    16'd63595: out <= 16'h01ED;
    16'd63596: out <= 16'hFF90;    16'd63597: out <= 16'hFFA2;    16'd63598: out <= 16'h0527;    16'd63599: out <= 16'hFA5F;
    16'd63600: out <= 16'hFF91;    16'd63601: out <= 16'hFC6A;    16'd63602: out <= 16'h0372;    16'd63603: out <= 16'hFE00;
    16'd63604: out <= 16'hFBCE;    16'd63605: out <= 16'hFC27;    16'd63606: out <= 16'h0208;    16'd63607: out <= 16'hFDEC;
    16'd63608: out <= 16'h0692;    16'd63609: out <= 16'h0302;    16'd63610: out <= 16'h0309;    16'd63611: out <= 16'hFD02;
    16'd63612: out <= 16'h02EF;    16'd63613: out <= 16'hFC3D;    16'd63614: out <= 16'h001A;    16'd63615: out <= 16'h0242;
    16'd63616: out <= 16'h0072;    16'd63617: out <= 16'h02E5;    16'd63618: out <= 16'hFBF6;    16'd63619: out <= 16'h0145;
    16'd63620: out <= 16'h0128;    16'd63621: out <= 16'hF9EC;    16'd63622: out <= 16'h00F1;    16'd63623: out <= 16'hFE04;
    16'd63624: out <= 16'hFF02;    16'd63625: out <= 16'hFA1F;    16'd63626: out <= 16'hFF9E;    16'd63627: out <= 16'h01C9;
    16'd63628: out <= 16'h002D;    16'd63629: out <= 16'hFC24;    16'd63630: out <= 16'h0117;    16'd63631: out <= 16'hFFC6;
    16'd63632: out <= 16'hFF3C;    16'd63633: out <= 16'hFE50;    16'd63634: out <= 16'hFFBC;    16'd63635: out <= 16'h0199;
    16'd63636: out <= 16'h013D;    16'd63637: out <= 16'hFD8F;    16'd63638: out <= 16'h00A2;    16'd63639: out <= 16'h076D;
    16'd63640: out <= 16'hFF53;    16'd63641: out <= 16'hFCBD;    16'd63642: out <= 16'h05B6;    16'd63643: out <= 16'hFD9A;
    16'd63644: out <= 16'h07DD;    16'd63645: out <= 16'h0143;    16'd63646: out <= 16'hFC1C;    16'd63647: out <= 16'h02A7;
    16'd63648: out <= 16'h0184;    16'd63649: out <= 16'h0001;    16'd63650: out <= 16'h0554;    16'd63651: out <= 16'h03AD;
    16'd63652: out <= 16'h063C;    16'd63653: out <= 16'hFFBF;    16'd63654: out <= 16'h0034;    16'd63655: out <= 16'h05EE;
    16'd63656: out <= 16'h047C;    16'd63657: out <= 16'h051C;    16'd63658: out <= 16'hFE81;    16'd63659: out <= 16'hFED2;
    16'd63660: out <= 16'hFB79;    16'd63661: out <= 16'h0984;    16'd63662: out <= 16'hFB55;    16'd63663: out <= 16'h03A6;
    16'd63664: out <= 16'h00A9;    16'd63665: out <= 16'hFFE0;    16'd63666: out <= 16'h091E;    16'd63667: out <= 16'h07C5;
    16'd63668: out <= 16'h00E6;    16'd63669: out <= 16'h0837;    16'd63670: out <= 16'h0336;    16'd63671: out <= 16'hFB23;
    16'd63672: out <= 16'hFE9C;    16'd63673: out <= 16'h05D1;    16'd63674: out <= 16'h071F;    16'd63675: out <= 16'h055D;
    16'd63676: out <= 16'h07D3;    16'd63677: out <= 16'h061C;    16'd63678: out <= 16'h0200;    16'd63679: out <= 16'h07C4;
    16'd63680: out <= 16'h0639;    16'd63681: out <= 16'h0908;    16'd63682: out <= 16'h0512;    16'd63683: out <= 16'h01F4;
    16'd63684: out <= 16'h0553;    16'd63685: out <= 16'h016D;    16'd63686: out <= 16'h0A8F;    16'd63687: out <= 16'h0265;
    16'd63688: out <= 16'hFC05;    16'd63689: out <= 16'hFE4B;    16'd63690: out <= 16'hFAD1;    16'd63691: out <= 16'hFE07;
    16'd63692: out <= 16'h02B2;    16'd63693: out <= 16'hFEC5;    16'd63694: out <= 16'hFE8C;    16'd63695: out <= 16'h02B1;
    16'd63696: out <= 16'h050B;    16'd63697: out <= 16'hFDED;    16'd63698: out <= 16'h0061;    16'd63699: out <= 16'h013F;
    16'd63700: out <= 16'h009A;    16'd63701: out <= 16'hFC3F;    16'd63702: out <= 16'h0178;    16'd63703: out <= 16'hF90A;
    16'd63704: out <= 16'hFB4A;    16'd63705: out <= 16'h0248;    16'd63706: out <= 16'h02CB;    16'd63707: out <= 16'hFBC9;
    16'd63708: out <= 16'h051A;    16'd63709: out <= 16'h019B;    16'd63710: out <= 16'h0153;    16'd63711: out <= 16'hFFB5;
    16'd63712: out <= 16'hFF06;    16'd63713: out <= 16'h0116;    16'd63714: out <= 16'hFC81;    16'd63715: out <= 16'hFFAC;
    16'd63716: out <= 16'hF9EE;    16'd63717: out <= 16'h065E;    16'd63718: out <= 16'h0243;    16'd63719: out <= 16'h022F;
    16'd63720: out <= 16'hFB03;    16'd63721: out <= 16'hFA85;    16'd63722: out <= 16'hFB90;    16'd63723: out <= 16'h03DF;
    16'd63724: out <= 16'h009C;    16'd63725: out <= 16'hFFC0;    16'd63726: out <= 16'h00BD;    16'd63727: out <= 16'h00D6;
    16'd63728: out <= 16'h04C1;    16'd63729: out <= 16'h00D8;    16'd63730: out <= 16'h003D;    16'd63731: out <= 16'hF8F2;
    16'd63732: out <= 16'h0265;    16'd63733: out <= 16'hFD6B;    16'd63734: out <= 16'hFCC8;    16'd63735: out <= 16'h03A1;
    16'd63736: out <= 16'h0236;    16'd63737: out <= 16'hFEA8;    16'd63738: out <= 16'hFFCE;    16'd63739: out <= 16'hF83E;
    16'd63740: out <= 16'h020C;    16'd63741: out <= 16'hFB29;    16'd63742: out <= 16'hF9F1;    16'd63743: out <= 16'hFE85;
    16'd63744: out <= 16'hFE0C;    16'd63745: out <= 16'h02AD;    16'd63746: out <= 16'h0009;    16'd63747: out <= 16'h02B8;
    16'd63748: out <= 16'hFDD3;    16'd63749: out <= 16'hFF04;    16'd63750: out <= 16'hFAB3;    16'd63751: out <= 16'hFFCF;
    16'd63752: out <= 16'h0067;    16'd63753: out <= 16'hFEF9;    16'd63754: out <= 16'h04CC;    16'd63755: out <= 16'hFFF5;
    16'd63756: out <= 16'h014F;    16'd63757: out <= 16'h0030;    16'd63758: out <= 16'h03D9;    16'd63759: out <= 16'h0138;
    16'd63760: out <= 16'hFC22;    16'd63761: out <= 16'hFACD;    16'd63762: out <= 16'hFAF4;    16'd63763: out <= 16'hFCEF;
    16'd63764: out <= 16'h0968;    16'd63765: out <= 16'h0905;    16'd63766: out <= 16'h0209;    16'd63767: out <= 16'hFB49;
    16'd63768: out <= 16'hFF76;    16'd63769: out <= 16'hF8D9;    16'd63770: out <= 16'h02AA;    16'd63771: out <= 16'hF767;
    16'd63772: out <= 16'h0C34;    16'd63773: out <= 16'hFA02;    16'd63774: out <= 16'hFCF3;    16'd63775: out <= 16'hF7E1;
    16'd63776: out <= 16'h0081;    16'd63777: out <= 16'hFE01;    16'd63778: out <= 16'h0375;    16'd63779: out <= 16'h0168;
    16'd63780: out <= 16'h0459;    16'd63781: out <= 16'h04D9;    16'd63782: out <= 16'h0213;    16'd63783: out <= 16'h0599;
    16'd63784: out <= 16'h06DF;    16'd63785: out <= 16'hFE40;    16'd63786: out <= 16'h04DA;    16'd63787: out <= 16'h00C9;
    16'd63788: out <= 16'h07B8;    16'd63789: out <= 16'h05DC;    16'd63790: out <= 16'h054D;    16'd63791: out <= 16'h08A9;
    16'd63792: out <= 16'h03E4;    16'd63793: out <= 16'h0B34;    16'd63794: out <= 16'h01A4;    16'd63795: out <= 16'h00F9;
    16'd63796: out <= 16'h063F;    16'd63797: out <= 16'h0503;    16'd63798: out <= 16'h00D0;    16'd63799: out <= 16'hFC11;
    16'd63800: out <= 16'hFF2E;    16'd63801: out <= 16'h01DA;    16'd63802: out <= 16'h0486;    16'd63803: out <= 16'h037A;
    16'd63804: out <= 16'h0685;    16'd63805: out <= 16'h04C1;    16'd63806: out <= 16'h01A0;    16'd63807: out <= 16'h075A;
    16'd63808: out <= 16'h0BBA;    16'd63809: out <= 16'h0088;    16'd63810: out <= 16'h04E5;    16'd63811: out <= 16'h015E;
    16'd63812: out <= 16'h0877;    16'd63813: out <= 16'h0301;    16'd63814: out <= 16'h00D4;    16'd63815: out <= 16'h03FC;
    16'd63816: out <= 16'h081F;    16'd63817: out <= 16'h0B5B;    16'd63818: out <= 16'hFEC5;    16'd63819: out <= 16'h0852;
    16'd63820: out <= 16'h02B6;    16'd63821: out <= 16'h05B4;    16'd63822: out <= 16'h0494;    16'd63823: out <= 16'h053B;
    16'd63824: out <= 16'h0224;    16'd63825: out <= 16'h0731;    16'd63826: out <= 16'h05E4;    16'd63827: out <= 16'h0214;
    16'd63828: out <= 16'h0851;    16'd63829: out <= 16'h0071;    16'd63830: out <= 16'h0608;    16'd63831: out <= 16'h05BB;
    16'd63832: out <= 16'h043B;    16'd63833: out <= 16'h0321;    16'd63834: out <= 16'hFFED;    16'd63835: out <= 16'h039F;
    16'd63836: out <= 16'h0C01;    16'd63837: out <= 16'h0431;    16'd63838: out <= 16'hFCCD;    16'd63839: out <= 16'h02B0;
    16'd63840: out <= 16'hFB6C;    16'd63841: out <= 16'h01E9;    16'd63842: out <= 16'h02DB;    16'd63843: out <= 16'h01B0;
    16'd63844: out <= 16'hFE0D;    16'd63845: out <= 16'h0030;    16'd63846: out <= 16'h02D3;    16'd63847: out <= 16'h026E;
    16'd63848: out <= 16'h007D;    16'd63849: out <= 16'hF889;    16'd63850: out <= 16'hFCBE;    16'd63851: out <= 16'h044A;
    16'd63852: out <= 16'hFF01;    16'd63853: out <= 16'h04D4;    16'd63854: out <= 16'h03CF;    16'd63855: out <= 16'hF846;
    16'd63856: out <= 16'h082C;    16'd63857: out <= 16'hFA07;    16'd63858: out <= 16'hFE1A;    16'd63859: out <= 16'hFD6D;
    16'd63860: out <= 16'h0318;    16'd63861: out <= 16'h0285;    16'd63862: out <= 16'h014C;    16'd63863: out <= 16'h03E5;
    16'd63864: out <= 16'hFF75;    16'd63865: out <= 16'hFC80;    16'd63866: out <= 16'hFFFB;    16'd63867: out <= 16'hFA7B;
    16'd63868: out <= 16'hFD6A;    16'd63869: out <= 16'hFFA3;    16'd63870: out <= 16'hFEC7;    16'd63871: out <= 16'hFF56;
    16'd63872: out <= 16'hFFED;    16'd63873: out <= 16'h08EE;    16'd63874: out <= 16'hFF8B;    16'd63875: out <= 16'h0601;
    16'd63876: out <= 16'h0197;    16'd63877: out <= 16'hFD7F;    16'd63878: out <= 16'h0100;    16'd63879: out <= 16'hFD94;
    16'd63880: out <= 16'hFACD;    16'd63881: out <= 16'hFEE0;    16'd63882: out <= 16'h00EF;    16'd63883: out <= 16'hF59B;
    16'd63884: out <= 16'hF652;    16'd63885: out <= 16'hFB96;    16'd63886: out <= 16'hF71A;    16'd63887: out <= 16'h00C1;
    16'd63888: out <= 16'h0209;    16'd63889: out <= 16'hF8A5;    16'd63890: out <= 16'h08B3;    16'd63891: out <= 16'hFFE9;
    16'd63892: out <= 16'hFAB8;    16'd63893: out <= 16'h03E6;    16'd63894: out <= 16'h02C6;    16'd63895: out <= 16'hFDC5;
    16'd63896: out <= 16'hFC4D;    16'd63897: out <= 16'hFD5C;    16'd63898: out <= 16'hFB61;    16'd63899: out <= 16'hFF4A;
    16'd63900: out <= 16'h000C;    16'd63901: out <= 16'h059D;    16'd63902: out <= 16'hFF43;    16'd63903: out <= 16'h03DB;
    16'd63904: out <= 16'h03A3;    16'd63905: out <= 16'h04FB;    16'd63906: out <= 16'h0043;    16'd63907: out <= 16'h0460;
    16'd63908: out <= 16'h02A6;    16'd63909: out <= 16'h00F9;    16'd63910: out <= 16'hFF16;    16'd63911: out <= 16'h0740;
    16'd63912: out <= 16'hFAC7;    16'd63913: out <= 16'hFEB5;    16'd63914: out <= 16'h0703;    16'd63915: out <= 16'h0C82;
    16'd63916: out <= 16'h054F;    16'd63917: out <= 16'h0634;    16'd63918: out <= 16'h04C1;    16'd63919: out <= 16'h01DD;
    16'd63920: out <= 16'hFEC4;    16'd63921: out <= 16'h0A96;    16'd63922: out <= 16'h03C9;    16'd63923: out <= 16'h0628;
    16'd63924: out <= 16'h009C;    16'd63925: out <= 16'h0748;    16'd63926: out <= 16'h022A;    16'd63927: out <= 16'hFFD6;
    16'd63928: out <= 16'h022C;    16'd63929: out <= 16'hFFE9;    16'd63930: out <= 16'h0252;    16'd63931: out <= 16'h0853;
    16'd63932: out <= 16'h00CF;    16'd63933: out <= 16'h00E4;    16'd63934: out <= 16'h0080;    16'd63935: out <= 16'hFD26;
    16'd63936: out <= 16'h0453;    16'd63937: out <= 16'hFDC7;    16'd63938: out <= 16'h0551;    16'd63939: out <= 16'h03B4;
    16'd63940: out <= 16'hFBE6;    16'd63941: out <= 16'hFF31;    16'd63942: out <= 16'hF277;    16'd63943: out <= 16'h0AB3;
    16'd63944: out <= 16'hFE73;    16'd63945: out <= 16'hFB31;    16'd63946: out <= 16'hF990;    16'd63947: out <= 16'hFBF3;
    16'd63948: out <= 16'hFCD5;    16'd63949: out <= 16'hF9CF;    16'd63950: out <= 16'h01D8;    16'd63951: out <= 16'hFDB9;
    16'd63952: out <= 16'hFFD2;    16'd63953: out <= 16'h01F4;    16'd63954: out <= 16'h0155;    16'd63955: out <= 16'h01FF;
    16'd63956: out <= 16'h02D4;    16'd63957: out <= 16'h034F;    16'd63958: out <= 16'h02F9;    16'd63959: out <= 16'hF878;
    16'd63960: out <= 16'h0027;    16'd63961: out <= 16'hFCF2;    16'd63962: out <= 16'hFA65;    16'd63963: out <= 16'hFC6D;
    16'd63964: out <= 16'h011A;    16'd63965: out <= 16'hFF66;    16'd63966: out <= 16'h0019;    16'd63967: out <= 16'h01AA;
    16'd63968: out <= 16'h06E0;    16'd63969: out <= 16'h0017;    16'd63970: out <= 16'hFF09;    16'd63971: out <= 16'hFDCC;
    16'd63972: out <= 16'hFF99;    16'd63973: out <= 16'hFEAF;    16'd63974: out <= 16'h02E6;    16'd63975: out <= 16'hFF07;
    16'd63976: out <= 16'hFCE1;    16'd63977: out <= 16'hFC51;    16'd63978: out <= 16'h0834;    16'd63979: out <= 16'h03E8;
    16'd63980: out <= 16'h04E3;    16'd63981: out <= 16'hF7C5;    16'd63982: out <= 16'h0368;    16'd63983: out <= 16'h0367;
    16'd63984: out <= 16'h002C;    16'd63985: out <= 16'h03C5;    16'd63986: out <= 16'hFFAA;    16'd63987: out <= 16'h06E3;
    16'd63988: out <= 16'hFCA1;    16'd63989: out <= 16'h01A0;    16'd63990: out <= 16'hFCF2;    16'd63991: out <= 16'hFC2F;
    16'd63992: out <= 16'h0324;    16'd63993: out <= 16'h0315;    16'd63994: out <= 16'hFD78;    16'd63995: out <= 16'h0509;
    16'd63996: out <= 16'h0232;    16'd63997: out <= 16'hFD4C;    16'd63998: out <= 16'hFA0B;    16'd63999: out <= 16'h0098;
    16'd64000: out <= 16'hFAEC;    16'd64001: out <= 16'h0482;    16'd64002: out <= 16'h03DC;    16'd64003: out <= 16'h0852;
    16'd64004: out <= 16'h0193;    16'd64005: out <= 16'hFFF8;    16'd64006: out <= 16'hFBBC;    16'd64007: out <= 16'hFBEC;
    16'd64008: out <= 16'hFE92;    16'd64009: out <= 16'h06C9;    16'd64010: out <= 16'h02B9;    16'd64011: out <= 16'h014C;
    16'd64012: out <= 16'hFE04;    16'd64013: out <= 16'h022B;    16'd64014: out <= 16'h02EA;    16'd64015: out <= 16'h0355;
    16'd64016: out <= 16'h01EF;    16'd64017: out <= 16'h0045;    16'd64018: out <= 16'hF82F;    16'd64019: out <= 16'hFDEA;
    16'd64020: out <= 16'hFFA5;    16'd64021: out <= 16'h048A;    16'd64022: out <= 16'hFEBF;    16'd64023: out <= 16'h034B;
    16'd64024: out <= 16'h0676;    16'd64025: out <= 16'h02BF;    16'd64026: out <= 16'hFDC4;    16'd64027: out <= 16'hFE0C;
    16'd64028: out <= 16'h0098;    16'd64029: out <= 16'h0475;    16'd64030: out <= 16'h0151;    16'd64031: out <= 16'hFB31;
    16'd64032: out <= 16'h013B;    16'd64033: out <= 16'h06AE;    16'd64034: out <= 16'h0810;    16'd64035: out <= 16'h043F;
    16'd64036: out <= 16'h02AB;    16'd64037: out <= 16'hF8FC;    16'd64038: out <= 16'hFDD9;    16'd64039: out <= 16'h0990;
    16'd64040: out <= 16'hFF19;    16'd64041: out <= 16'hFC07;    16'd64042: out <= 16'h069E;    16'd64043: out <= 16'h04E1;
    16'd64044: out <= 16'h0615;    16'd64045: out <= 16'h0976;    16'd64046: out <= 16'h0630;    16'd64047: out <= 16'h028F;
    16'd64048: out <= 16'hFF88;    16'd64049: out <= 16'hFF80;    16'd64050: out <= 16'h0722;    16'd64051: out <= 16'h037C;
    16'd64052: out <= 16'h0B01;    16'd64053: out <= 16'h0424;    16'd64054: out <= 16'hFE31;    16'd64055: out <= 16'h0426;
    16'd64056: out <= 16'h0568;    16'd64057: out <= 16'h06E4;    16'd64058: out <= 16'h0092;    16'd64059: out <= 16'h02DC;
    16'd64060: out <= 16'h052C;    16'd64061: out <= 16'h0F6E;    16'd64062: out <= 16'hFA5C;    16'd64063: out <= 16'h04EC;
    16'd64064: out <= 16'h08DB;    16'd64065: out <= 16'h0181;    16'd64066: out <= 16'hFDB6;    16'd64067: out <= 16'h005D;
    16'd64068: out <= 16'h0783;    16'd64069: out <= 16'h0259;    16'd64070: out <= 16'h0256;    16'd64071: out <= 16'h07FC;
    16'd64072: out <= 16'h0980;    16'd64073: out <= 16'h04D6;    16'd64074: out <= 16'hFE71;    16'd64075: out <= 16'hFB70;
    16'd64076: out <= 16'h0B34;    16'd64077: out <= 16'h06FA;    16'd64078: out <= 16'hFCA6;    16'd64079: out <= 16'h0553;
    16'd64080: out <= 16'h0282;    16'd64081: out <= 16'hFEFA;    16'd64082: out <= 16'h02BA;    16'd64083: out <= 16'h068D;
    16'd64084: out <= 16'h0018;    16'd64085: out <= 16'h02C2;    16'd64086: out <= 16'h097F;    16'd64087: out <= 16'h0A03;
    16'd64088: out <= 16'h0BE9;    16'd64089: out <= 16'h010B;    16'd64090: out <= 16'h06E2;    16'd64091: out <= 16'h0509;
    16'd64092: out <= 16'hFE0B;    16'd64093: out <= 16'hFF75;    16'd64094: out <= 16'hFD52;    16'd64095: out <= 16'hFD8B;
    16'd64096: out <= 16'h0222;    16'd64097: out <= 16'h036F;    16'd64098: out <= 16'h00C5;    16'd64099: out <= 16'hF922;
    16'd64100: out <= 16'h01E8;    16'd64101: out <= 16'hFDE2;    16'd64102: out <= 16'hFB56;    16'd64103: out <= 16'h0231;
    16'd64104: out <= 16'h0307;    16'd64105: out <= 16'h0489;    16'd64106: out <= 16'h079B;    16'd64107: out <= 16'h0C07;
    16'd64108: out <= 16'hFE96;    16'd64109: out <= 16'h01E5;    16'd64110: out <= 16'h03D3;    16'd64111: out <= 16'hFC05;
    16'd64112: out <= 16'h039F;    16'd64113: out <= 16'h005A;    16'd64114: out <= 16'hF670;    16'd64115: out <= 16'h006D;
    16'd64116: out <= 16'hFCC5;    16'd64117: out <= 16'hFBA2;    16'd64118: out <= 16'h05A2;    16'd64119: out <= 16'hFDCC;
    16'd64120: out <= 16'hF790;    16'd64121: out <= 16'hF5E0;    16'd64122: out <= 16'h04BA;    16'd64123: out <= 16'hFDEF;
    16'd64124: out <= 16'hFB0C;    16'd64125: out <= 16'h0433;    16'd64126: out <= 16'hFF5A;    16'd64127: out <= 16'hFBB8;
    16'd64128: out <= 16'hFEF4;    16'd64129: out <= 16'hF8B4;    16'd64130: out <= 16'hFEA9;    16'd64131: out <= 16'hFEAC;
    16'd64132: out <= 16'hFE11;    16'd64133: out <= 16'hFEDC;    16'd64134: out <= 16'h009D;    16'd64135: out <= 16'hFAAC;
    16'd64136: out <= 16'h03A8;    16'd64137: out <= 16'hFCD4;    16'd64138: out <= 16'hF820;    16'd64139: out <= 16'h08AE;
    16'd64140: out <= 16'h07A0;    16'd64141: out <= 16'hFFBA;    16'd64142: out <= 16'h02D4;    16'd64143: out <= 16'hFF98;
    16'd64144: out <= 16'hF633;    16'd64145: out <= 16'hFECF;    16'd64146: out <= 16'hF4FF;    16'd64147: out <= 16'h07D3;
    16'd64148: out <= 16'hFDDE;    16'd64149: out <= 16'h0360;    16'd64150: out <= 16'hFF1B;    16'd64151: out <= 16'hFFB7;
    16'd64152: out <= 16'hFF65;    16'd64153: out <= 16'h0387;    16'd64154: out <= 16'h0637;    16'd64155: out <= 16'h08AB;
    16'd64156: out <= 16'h00FE;    16'd64157: out <= 16'h0680;    16'd64158: out <= 16'h05EF;    16'd64159: out <= 16'h01D8;
    16'd64160: out <= 16'h0103;    16'd64161: out <= 16'h0296;    16'd64162: out <= 16'h0789;    16'd64163: out <= 16'h027B;
    16'd64164: out <= 16'hFF18;    16'd64165: out <= 16'h0705;    16'd64166: out <= 16'h03EE;    16'd64167: out <= 16'h09F6;
    16'd64168: out <= 16'h0401;    16'd64169: out <= 16'h0209;    16'd64170: out <= 16'h019E;    16'd64171: out <= 16'h0751;
    16'd64172: out <= 16'h03F7;    16'd64173: out <= 16'hFFE7;    16'd64174: out <= 16'hFB51;    16'd64175: out <= 16'h0732;
    16'd64176: out <= 16'h0510;    16'd64177: out <= 16'h04C3;    16'd64178: out <= 16'h01A9;    16'd64179: out <= 16'h099E;
    16'd64180: out <= 16'h0502;    16'd64181: out <= 16'h03C1;    16'd64182: out <= 16'h05DE;    16'd64183: out <= 16'hFF10;
    16'd64184: out <= 16'h01E9;    16'd64185: out <= 16'h04D8;    16'd64186: out <= 16'h01C8;    16'd64187: out <= 16'h0647;
    16'd64188: out <= 16'h04EA;    16'd64189: out <= 16'hFDFC;    16'd64190: out <= 16'h04C5;    16'd64191: out <= 16'h02AA;
    16'd64192: out <= 16'h0A2F;    16'd64193: out <= 16'hFFD9;    16'd64194: out <= 16'h0867;    16'd64195: out <= 16'h06BB;
    16'd64196: out <= 16'h0559;    16'd64197: out <= 16'h0000;    16'd64198: out <= 16'hFAD9;    16'd64199: out <= 16'h0613;
    16'd64200: out <= 16'hFB23;    16'd64201: out <= 16'h004C;    16'd64202: out <= 16'h0131;    16'd64203: out <= 16'hFEDC;
    16'd64204: out <= 16'hFCC8;    16'd64205: out <= 16'h0655;    16'd64206: out <= 16'h07AE;    16'd64207: out <= 16'h03CB;
    16'd64208: out <= 16'h0438;    16'd64209: out <= 16'hFC7C;    16'd64210: out <= 16'hFDC5;    16'd64211: out <= 16'h02E9;
    16'd64212: out <= 16'h008C;    16'd64213: out <= 16'hFDE5;    16'd64214: out <= 16'h0040;    16'd64215: out <= 16'hFE3D;
    16'd64216: out <= 16'h010E;    16'd64217: out <= 16'h047A;    16'd64218: out <= 16'hFE92;    16'd64219: out <= 16'h02D4;
    16'd64220: out <= 16'hFFBB;    16'd64221: out <= 16'hFD8C;    16'd64222: out <= 16'h0162;    16'd64223: out <= 16'h04B1;
    16'd64224: out <= 16'h020A;    16'd64225: out <= 16'h038B;    16'd64226: out <= 16'h00BC;    16'd64227: out <= 16'h00F8;
    16'd64228: out <= 16'h065D;    16'd64229: out <= 16'hFDCE;    16'd64230: out <= 16'h027D;    16'd64231: out <= 16'h0704;
    16'd64232: out <= 16'hFBBA;    16'd64233: out <= 16'hFE07;    16'd64234: out <= 16'h0028;    16'd64235: out <= 16'h0319;
    16'd64236: out <= 16'hF9CE;    16'd64237: out <= 16'h05DC;    16'd64238: out <= 16'h045D;    16'd64239: out <= 16'hFFCE;
    16'd64240: out <= 16'hFAAF;    16'd64241: out <= 16'h015F;    16'd64242: out <= 16'hFE30;    16'd64243: out <= 16'hFC76;
    16'd64244: out <= 16'hFFD5;    16'd64245: out <= 16'hFB03;    16'd64246: out <= 16'hF9DF;    16'd64247: out <= 16'hFB72;
    16'd64248: out <= 16'hFA07;    16'd64249: out <= 16'hFFB5;    16'd64250: out <= 16'h034A;    16'd64251: out <= 16'h03E8;
    16'd64252: out <= 16'hFC68;    16'd64253: out <= 16'h025C;    16'd64254: out <= 16'hFDDE;    16'd64255: out <= 16'hFF13;
    16'd64256: out <= 16'hFFE4;    16'd64257: out <= 16'h00A3;    16'd64258: out <= 16'hFFB4;    16'd64259: out <= 16'hFEDD;
    16'd64260: out <= 16'h0180;    16'd64261: out <= 16'hFA08;    16'd64262: out <= 16'h03A0;    16'd64263: out <= 16'hFD1F;
    16'd64264: out <= 16'hFC55;    16'd64265: out <= 16'hFC35;    16'd64266: out <= 16'h06EF;    16'd64267: out <= 16'h071B;
    16'd64268: out <= 16'hFA1B;    16'd64269: out <= 16'hF938;    16'd64270: out <= 16'h01A8;    16'd64271: out <= 16'h03BB;
    16'd64272: out <= 16'h057A;    16'd64273: out <= 16'h0268;    16'd64274: out <= 16'hFCBD;    16'd64275: out <= 16'h01E4;
    16'd64276: out <= 16'hFC93;    16'd64277: out <= 16'h0864;    16'd64278: out <= 16'h081A;    16'd64279: out <= 16'h014E;
    16'd64280: out <= 16'hFABE;    16'd64281: out <= 16'hFDEA;    16'd64282: out <= 16'h0264;    16'd64283: out <= 16'h0939;
    16'd64284: out <= 16'hFFAA;    16'd64285: out <= 16'hFAF4;    16'd64286: out <= 16'h0093;    16'd64287: out <= 16'hFF98;
    16'd64288: out <= 16'hFAD6;    16'd64289: out <= 16'h03D4;    16'd64290: out <= 16'hF7E6;    16'd64291: out <= 16'hFE64;
    16'd64292: out <= 16'h039C;    16'd64293: out <= 16'hFF79;    16'd64294: out <= 16'h02CC;    16'd64295: out <= 16'hFDD2;
    16'd64296: out <= 16'h0094;    16'd64297: out <= 16'h0683;    16'd64298: out <= 16'h036E;    16'd64299: out <= 16'h00B9;
    16'd64300: out <= 16'h085A;    16'd64301: out <= 16'hFE94;    16'd64302: out <= 16'h0206;    16'd64303: out <= 16'h0AFB;
    16'd64304: out <= 16'h0098;    16'd64305: out <= 16'h0939;    16'd64306: out <= 16'hFECF;    16'd64307: out <= 16'h0A75;
    16'd64308: out <= 16'h017E;    16'd64309: out <= 16'hFA21;    16'd64310: out <= 16'h05B7;    16'd64311: out <= 16'hFF95;
    16'd64312: out <= 16'h0D27;    16'd64313: out <= 16'hFC83;    16'd64314: out <= 16'h057B;    16'd64315: out <= 16'h050D;
    16'd64316: out <= 16'h0662;    16'd64317: out <= 16'h0385;    16'd64318: out <= 16'h07DA;    16'd64319: out <= 16'hFFFA;
    16'd64320: out <= 16'h08F9;    16'd64321: out <= 16'h02E1;    16'd64322: out <= 16'h0455;    16'd64323: out <= 16'h046E;
    16'd64324: out <= 16'h07AD;    16'd64325: out <= 16'h0238;    16'd64326: out <= 16'h0340;    16'd64327: out <= 16'h04AA;
    16'd64328: out <= 16'h05DE;    16'd64329: out <= 16'h01EB;    16'd64330: out <= 16'h0933;    16'd64331: out <= 16'h03F3;
    16'd64332: out <= 16'h0981;    16'd64333: out <= 16'h03BB;    16'd64334: out <= 16'h0348;    16'd64335: out <= 16'h0A50;
    16'd64336: out <= 16'h0289;    16'd64337: out <= 16'hFE6A;    16'd64338: out <= 16'h06CD;    16'd64339: out <= 16'h0570;
    16'd64340: out <= 16'h0222;    16'd64341: out <= 16'h0319;    16'd64342: out <= 16'h0CBC;    16'd64343: out <= 16'h0528;
    16'd64344: out <= 16'h03EA;    16'd64345: out <= 16'h0101;    16'd64346: out <= 16'h01CE;    16'd64347: out <= 16'h06B3;
    16'd64348: out <= 16'h09AD;    16'd64349: out <= 16'hFB45;    16'd64350: out <= 16'h010B;    16'd64351: out <= 16'hFFC7;
    16'd64352: out <= 16'h03E0;    16'd64353: out <= 16'hFF06;    16'd64354: out <= 16'hFCF2;    16'd64355: out <= 16'h014E;
    16'd64356: out <= 16'hFC98;    16'd64357: out <= 16'hFF58;    16'd64358: out <= 16'hFEA9;    16'd64359: out <= 16'h03E7;
    16'd64360: out <= 16'hFEBC;    16'd64361: out <= 16'h038E;    16'd64362: out <= 16'h03CC;    16'd64363: out <= 16'h0158;
    16'd64364: out <= 16'h026C;    16'd64365: out <= 16'hFC40;    16'd64366: out <= 16'hFD95;    16'd64367: out <= 16'h040D;
    16'd64368: out <= 16'h00E3;    16'd64369: out <= 16'hFEA5;    16'd64370: out <= 16'h005E;    16'd64371: out <= 16'h0494;
    16'd64372: out <= 16'hFD4A;    16'd64373: out <= 16'h013A;    16'd64374: out <= 16'h0374;    16'd64375: out <= 16'h0323;
    16'd64376: out <= 16'h00E6;    16'd64377: out <= 16'hFCB7;    16'd64378: out <= 16'h0359;    16'd64379: out <= 16'h02B3;
    16'd64380: out <= 16'hFC90;    16'd64381: out <= 16'h01FA;    16'd64382: out <= 16'h0356;    16'd64383: out <= 16'hFFEC;
    16'd64384: out <= 16'hF914;    16'd64385: out <= 16'h06C4;    16'd64386: out <= 16'hFFED;    16'd64387: out <= 16'h00B4;
    16'd64388: out <= 16'hFD95;    16'd64389: out <= 16'hFB9F;    16'd64390: out <= 16'hFCD2;    16'd64391: out <= 16'hFA1F;
    16'd64392: out <= 16'h0869;    16'd64393: out <= 16'hFD95;    16'd64394: out <= 16'h0463;    16'd64395: out <= 16'hF810;
    16'd64396: out <= 16'h008C;    16'd64397: out <= 16'h0043;    16'd64398: out <= 16'h0658;    16'd64399: out <= 16'hFF01;
    16'd64400: out <= 16'h04CA;    16'd64401: out <= 16'hFEF2;    16'd64402: out <= 16'hFF76;    16'd64403: out <= 16'hFCD8;
    16'd64404: out <= 16'h097F;    16'd64405: out <= 16'h00FC;    16'd64406: out <= 16'hFCA4;    16'd64407: out <= 16'h01C8;
    16'd64408: out <= 16'h00F7;    16'd64409: out <= 16'hFC7E;    16'd64410: out <= 16'h0231;    16'd64411: out <= 16'hFD4A;
    16'd64412: out <= 16'hF987;    16'd64413: out <= 16'hFC9A;    16'd64414: out <= 16'hFB04;    16'd64415: out <= 16'hFDA2;
    16'd64416: out <= 16'h03FD;    16'd64417: out <= 16'hFD83;    16'd64418: out <= 16'h004A;    16'd64419: out <= 16'hFFD6;
    16'd64420: out <= 16'h0854;    16'd64421: out <= 16'h0756;    16'd64422: out <= 16'h04D5;    16'd64423: out <= 16'h049A;
    16'd64424: out <= 16'h057F;    16'd64425: out <= 16'h0635;    16'd64426: out <= 16'h056F;    16'd64427: out <= 16'h0065;
    16'd64428: out <= 16'h08D3;    16'd64429: out <= 16'h01E4;    16'd64430: out <= 16'hFFE1;    16'd64431: out <= 16'h0691;
    16'd64432: out <= 16'hFB4E;    16'd64433: out <= 16'h047F;    16'd64434: out <= 16'h0562;    16'd64435: out <= 16'hFEBC;
    16'd64436: out <= 16'h066E;    16'd64437: out <= 16'hFB18;    16'd64438: out <= 16'h05A2;    16'd64439: out <= 16'h02BE;
    16'd64440: out <= 16'hFF41;    16'd64441: out <= 16'h0FFF;    16'd64442: out <= 16'h04F1;    16'd64443: out <= 16'h0039;
    16'd64444: out <= 16'h07A1;    16'd64445: out <= 16'h05DF;    16'd64446: out <= 16'h04BC;    16'd64447: out <= 16'h05E2;
    16'd64448: out <= 16'h0718;    16'd64449: out <= 16'h01C3;    16'd64450: out <= 16'hFF7E;    16'd64451: out <= 16'h0677;
    16'd64452: out <= 16'h050C;    16'd64453: out <= 16'hFE65;    16'd64454: out <= 16'h0692;    16'd64455: out <= 16'hFCCF;
    16'd64456: out <= 16'h0214;    16'd64457: out <= 16'h0440;    16'd64458: out <= 16'h0566;    16'd64459: out <= 16'hFC30;
    16'd64460: out <= 16'h0164;    16'd64461: out <= 16'h0278;    16'd64462: out <= 16'hFEB0;    16'd64463: out <= 16'hFCD7;
    16'd64464: out <= 16'h01AB;    16'd64465: out <= 16'hFECA;    16'd64466: out <= 16'h03AE;    16'd64467: out <= 16'h0453;
    16'd64468: out <= 16'hFE1C;    16'd64469: out <= 16'h017D;    16'd64470: out <= 16'hF946;    16'd64471: out <= 16'h0255;
    16'd64472: out <= 16'h0084;    16'd64473: out <= 16'h000C;    16'd64474: out <= 16'h0033;    16'd64475: out <= 16'hF8EF;
    16'd64476: out <= 16'h0183;    16'd64477: out <= 16'h022E;    16'd64478: out <= 16'hFB39;    16'd64479: out <= 16'h015C;
    16'd64480: out <= 16'h00DC;    16'd64481: out <= 16'hFE11;    16'd64482: out <= 16'h0511;    16'd64483: out <= 16'h054D;
    16'd64484: out <= 16'h0090;    16'd64485: out <= 16'hFDD2;    16'd64486: out <= 16'hFCFF;    16'd64487: out <= 16'h0111;
    16'd64488: out <= 16'h0000;    16'd64489: out <= 16'h01C2;    16'd64490: out <= 16'h04CD;    16'd64491: out <= 16'hF91E;
    16'd64492: out <= 16'hFF6C;    16'd64493: out <= 16'hFDDB;    16'd64494: out <= 16'h00DB;    16'd64495: out <= 16'hFB8D;
    16'd64496: out <= 16'h01B1;    16'd64497: out <= 16'h070C;    16'd64498: out <= 16'hFD9C;    16'd64499: out <= 16'h00AF;
    16'd64500: out <= 16'hFFE0;    16'd64501: out <= 16'h0371;    16'd64502: out <= 16'hFD73;    16'd64503: out <= 16'hFD1A;
    16'd64504: out <= 16'hFD46;    16'd64505: out <= 16'h053E;    16'd64506: out <= 16'hFADA;    16'd64507: out <= 16'h069D;
    16'd64508: out <= 16'hFFD3;    16'd64509: out <= 16'hFF3B;    16'd64510: out <= 16'hFD60;    16'd64511: out <= 16'hFF82;
    16'd64512: out <= 16'h05AC;    16'd64513: out <= 16'hFDB7;    16'd64514: out <= 16'h011F;    16'd64515: out <= 16'h0729;
    16'd64516: out <= 16'h0806;    16'd64517: out <= 16'h03B3;    16'd64518: out <= 16'h0021;    16'd64519: out <= 16'hFCB5;
    16'd64520: out <= 16'hFE6F;    16'd64521: out <= 16'h009D;    16'd64522: out <= 16'hFC00;    16'd64523: out <= 16'hFF25;
    16'd64524: out <= 16'h01EF;    16'd64525: out <= 16'hFD7D;    16'd64526: out <= 16'hFB79;    16'd64527: out <= 16'hFCC9;
    16'd64528: out <= 16'h009F;    16'd64529: out <= 16'h04B9;    16'd64530: out <= 16'hFED3;    16'd64531: out <= 16'h01B4;
    16'd64532: out <= 16'hFEC1;    16'd64533: out <= 16'hFCF6;    16'd64534: out <= 16'h03A3;    16'd64535: out <= 16'h0127;
    16'd64536: out <= 16'hFB56;    16'd64537: out <= 16'hF7C5;    16'd64538: out <= 16'h053E;    16'd64539: out <= 16'hFFF7;
    16'd64540: out <= 16'h0109;    16'd64541: out <= 16'hF7BC;    16'd64542: out <= 16'h02B6;    16'd64543: out <= 16'h0333;
    16'd64544: out <= 16'h01BA;    16'd64545: out <= 16'h08EA;    16'd64546: out <= 16'h00E8;    16'd64547: out <= 16'h0DE8;
    16'd64548: out <= 16'h0564;    16'd64549: out <= 16'h0168;    16'd64550: out <= 16'h0549;    16'd64551: out <= 16'h0A8D;
    16'd64552: out <= 16'h01C4;    16'd64553: out <= 16'hFDBA;    16'd64554: out <= 16'hFE24;    16'd64555: out <= 16'h0B65;
    16'd64556: out <= 16'h0237;    16'd64557: out <= 16'h000F;    16'd64558: out <= 16'h0298;    16'd64559: out <= 16'h003B;
    16'd64560: out <= 16'h0415;    16'd64561: out <= 16'hFF5E;    16'd64562: out <= 16'h085B;    16'd64563: out <= 16'h086D;
    16'd64564: out <= 16'hFE00;    16'd64565: out <= 16'h046D;    16'd64566: out <= 16'h020A;    16'd64567: out <= 16'h065F;
    16'd64568: out <= 16'hFCDA;    16'd64569: out <= 16'h01EC;    16'd64570: out <= 16'h003E;    16'd64571: out <= 16'h0ADB;
    16'd64572: out <= 16'h044F;    16'd64573: out <= 16'h020C;    16'd64574: out <= 16'h04F2;    16'd64575: out <= 16'h0519;
    16'd64576: out <= 16'h05E1;    16'd64577: out <= 16'hFDAB;    16'd64578: out <= 16'h043B;    16'd64579: out <= 16'h06FF;
    16'd64580: out <= 16'h0870;    16'd64581: out <= 16'h0606;    16'd64582: out <= 16'h07C0;    16'd64583: out <= 16'h0716;
    16'd64584: out <= 16'h08E7;    16'd64585: out <= 16'h0586;    16'd64586: out <= 16'h0694;    16'd64587: out <= 16'h0793;
    16'd64588: out <= 16'h0248;    16'd64589: out <= 16'h019C;    16'd64590: out <= 16'hFF67;    16'd64591: out <= 16'hFCBF;
    16'd64592: out <= 16'h0499;    16'd64593: out <= 16'h08BC;    16'd64594: out <= 16'hFEAA;    16'd64595: out <= 16'h035D;
    16'd64596: out <= 16'h017F;    16'd64597: out <= 16'h036F;    16'd64598: out <= 16'h084B;    16'd64599: out <= 16'h0B6C;
    16'd64600: out <= 16'h03DA;    16'd64601: out <= 16'h03E4;    16'd64602: out <= 16'h017D;    16'd64603: out <= 16'h00DE;
    16'd64604: out <= 16'hFD5C;    16'd64605: out <= 16'h0284;    16'd64606: out <= 16'hF607;    16'd64607: out <= 16'h01F9;
    16'd64608: out <= 16'h0066;    16'd64609: out <= 16'h01DA;    16'd64610: out <= 16'h0187;    16'd64611: out <= 16'h04A9;
    16'd64612: out <= 16'h05C9;    16'd64613: out <= 16'h04DB;    16'd64614: out <= 16'h060E;    16'd64615: out <= 16'h04C1;
    16'd64616: out <= 16'h01BC;    16'd64617: out <= 16'h02D1;    16'd64618: out <= 16'hFC0F;    16'd64619: out <= 16'h01C1;
    16'd64620: out <= 16'h000D;    16'd64621: out <= 16'h0180;    16'd64622: out <= 16'hFEBC;    16'd64623: out <= 16'h039C;
    16'd64624: out <= 16'h04D9;    16'd64625: out <= 16'hFAB9;    16'd64626: out <= 16'h013A;    16'd64627: out <= 16'h0DCC;
    16'd64628: out <= 16'h0185;    16'd64629: out <= 16'hFE52;    16'd64630: out <= 16'h06E0;    16'd64631: out <= 16'h052C;
    16'd64632: out <= 16'h07B6;    16'd64633: out <= 16'h02A0;    16'd64634: out <= 16'hFFB3;    16'd64635: out <= 16'hFE7C;
    16'd64636: out <= 16'h05B1;    16'd64637: out <= 16'h04A2;    16'd64638: out <= 16'h0126;    16'd64639: out <= 16'h0013;
    16'd64640: out <= 16'hFDE7;    16'd64641: out <= 16'hFDA2;    16'd64642: out <= 16'h0206;    16'd64643: out <= 16'hFF25;
    16'd64644: out <= 16'hFF19;    16'd64645: out <= 16'h023B;    16'd64646: out <= 16'h03EF;    16'd64647: out <= 16'hF839;
    16'd64648: out <= 16'hFC84;    16'd64649: out <= 16'hF5B7;    16'd64650: out <= 16'h07B4;    16'd64651: out <= 16'h010E;
    16'd64652: out <= 16'h016D;    16'd64653: out <= 16'hFA80;    16'd64654: out <= 16'hF95F;    16'd64655: out <= 16'h01DE;
    16'd64656: out <= 16'h04FD;    16'd64657: out <= 16'hFAB0;    16'd64658: out <= 16'h0216;    16'd64659: out <= 16'hFB2B;
    16'd64660: out <= 16'h0010;    16'd64661: out <= 16'h023C;    16'd64662: out <= 16'hFE97;    16'd64663: out <= 16'hFE87;
    16'd64664: out <= 16'h04B3;    16'd64665: out <= 16'h0121;    16'd64666: out <= 16'h04DE;    16'd64667: out <= 16'h0276;
    16'd64668: out <= 16'hF873;    16'd64669: out <= 16'hF9BF;    16'd64670: out <= 16'h003B;    16'd64671: out <= 16'h0BE3;
    16'd64672: out <= 16'h061D;    16'd64673: out <= 16'hFB0B;    16'd64674: out <= 16'hFECD;    16'd64675: out <= 16'hFDCF;
    16'd64676: out <= 16'h01B1;    16'd64677: out <= 16'h0115;    16'd64678: out <= 16'h0856;    16'd64679: out <= 16'h00CB;
    16'd64680: out <= 16'h0890;    16'd64681: out <= 16'h0350;    16'd64682: out <= 16'hFEF5;    16'd64683: out <= 16'h0293;
    16'd64684: out <= 16'h026F;    16'd64685: out <= 16'h033A;    16'd64686: out <= 16'h01DF;    16'd64687: out <= 16'h092D;
    16'd64688: out <= 16'h08BE;    16'd64689: out <= 16'h0445;    16'd64690: out <= 16'h0A48;    16'd64691: out <= 16'h046F;
    16'd64692: out <= 16'h0223;    16'd64693: out <= 16'h01B1;    16'd64694: out <= 16'h04F5;    16'd64695: out <= 16'h038C;
    16'd64696: out <= 16'h0407;    16'd64697: out <= 16'h02BE;    16'd64698: out <= 16'h1108;    16'd64699: out <= 16'h04D9;
    16'd64700: out <= 16'hFF7E;    16'd64701: out <= 16'h058B;    16'd64702: out <= 16'h01F8;    16'd64703: out <= 16'hFF97;
    16'd64704: out <= 16'hFDFB;    16'd64705: out <= 16'h05C6;    16'd64706: out <= 16'h0896;    16'd64707: out <= 16'h0B4E;
    16'd64708: out <= 16'h03F0;    16'd64709: out <= 16'hFEED;    16'd64710: out <= 16'hFEE3;    16'd64711: out <= 16'hF8BE;
    16'd64712: out <= 16'h01EE;    16'd64713: out <= 16'hFA34;    16'd64714: out <= 16'h0169;    16'd64715: out <= 16'hFECC;
    16'd64716: out <= 16'h016A;    16'd64717: out <= 16'h0442;    16'd64718: out <= 16'h0390;    16'd64719: out <= 16'h0421;
    16'd64720: out <= 16'h0165;    16'd64721: out <= 16'h05A6;    16'd64722: out <= 16'h0878;    16'd64723: out <= 16'hFD4A;
    16'd64724: out <= 16'hF5DC;    16'd64725: out <= 16'h013C;    16'd64726: out <= 16'hFA56;    16'd64727: out <= 16'hF577;
    16'd64728: out <= 16'hFBF2;    16'd64729: out <= 16'h01F3;    16'd64730: out <= 16'h00D4;    16'd64731: out <= 16'hFD34;
    16'd64732: out <= 16'h0092;    16'd64733: out <= 16'hFFAC;    16'd64734: out <= 16'hFFBD;    16'd64735: out <= 16'h01A8;
    16'd64736: out <= 16'hFD37;    16'd64737: out <= 16'h02B3;    16'd64738: out <= 16'h0245;    16'd64739: out <= 16'h0351;
    16'd64740: out <= 16'h0049;    16'd64741: out <= 16'h002D;    16'd64742: out <= 16'h024A;    16'd64743: out <= 16'h0243;
    16'd64744: out <= 16'hFC2E;    16'd64745: out <= 16'hFF4A;    16'd64746: out <= 16'hFC6E;    16'd64747: out <= 16'hFE7A;
    16'd64748: out <= 16'hF80A;    16'd64749: out <= 16'h04EB;    16'd64750: out <= 16'hFF42;    16'd64751: out <= 16'h0122;
    16'd64752: out <= 16'hFFD2;    16'd64753: out <= 16'h0448;    16'd64754: out <= 16'h01E5;    16'd64755: out <= 16'hFD95;
    16'd64756: out <= 16'h0118;    16'd64757: out <= 16'hFD76;    16'd64758: out <= 16'hFE47;    16'd64759: out <= 16'hFE78;
    16'd64760: out <= 16'hFFBA;    16'd64761: out <= 16'hFE1E;    16'd64762: out <= 16'hFACC;    16'd64763: out <= 16'h0139;
    16'd64764: out <= 16'hFFE0;    16'd64765: out <= 16'hF8C4;    16'd64766: out <= 16'hFF83;    16'd64767: out <= 16'hFDF6;
    16'd64768: out <= 16'h0507;    16'd64769: out <= 16'hFC00;    16'd64770: out <= 16'h0124;    16'd64771: out <= 16'hFD00;
    16'd64772: out <= 16'h00FC;    16'd64773: out <= 16'hFF2C;    16'd64774: out <= 16'hFC67;    16'd64775: out <= 16'h07D8;
    16'd64776: out <= 16'h0545;    16'd64777: out <= 16'h0414;    16'd64778: out <= 16'h055E;    16'd64779: out <= 16'hFFE7;
    16'd64780: out <= 16'hFE09;    16'd64781: out <= 16'h05E6;    16'd64782: out <= 16'h0571;    16'd64783: out <= 16'h053B;
    16'd64784: out <= 16'hF95C;    16'd64785: out <= 16'h05C1;    16'd64786: out <= 16'hFDA0;    16'd64787: out <= 16'hFC23;
    16'd64788: out <= 16'h0809;    16'd64789: out <= 16'h0063;    16'd64790: out <= 16'h0043;    16'd64791: out <= 16'h00F7;
    16'd64792: out <= 16'h0155;    16'd64793: out <= 16'hFFFF;    16'd64794: out <= 16'h01D3;    16'd64795: out <= 16'hFEE4;
    16'd64796: out <= 16'h030A;    16'd64797: out <= 16'hFFD9;    16'd64798: out <= 16'hFD5A;    16'd64799: out <= 16'h019F;
    16'd64800: out <= 16'h0547;    16'd64801: out <= 16'hFBD4;    16'd64802: out <= 16'h05BB;    16'd64803: out <= 16'h04BD;
    16'd64804: out <= 16'h067E;    16'd64805: out <= 16'h00D8;    16'd64806: out <= 16'h06AC;    16'd64807: out <= 16'h053E;
    16'd64808: out <= 16'h0475;    16'd64809: out <= 16'h0D81;    16'd64810: out <= 16'hFEBA;    16'd64811: out <= 16'h089D;
    16'd64812: out <= 16'h0819;    16'd64813: out <= 16'h0811;    16'd64814: out <= 16'h073A;    16'd64815: out <= 16'h06EF;
    16'd64816: out <= 16'h01E7;    16'd64817: out <= 16'h00B5;    16'd64818: out <= 16'h040F;    16'd64819: out <= 16'h03FD;
    16'd64820: out <= 16'h053F;    16'd64821: out <= 16'hFF7D;    16'd64822: out <= 16'h0822;    16'd64823: out <= 16'h085D;
    16'd64824: out <= 16'h0144;    16'd64825: out <= 16'h0121;    16'd64826: out <= 16'h0507;    16'd64827: out <= 16'h03E0;
    16'd64828: out <= 16'h0236;    16'd64829: out <= 16'h00F9;    16'd64830: out <= 16'h0254;    16'd64831: out <= 16'h03B2;
    16'd64832: out <= 16'h0112;    16'd64833: out <= 16'hFF42;    16'd64834: out <= 16'h04F1;    16'd64835: out <= 16'h01C5;
    16'd64836: out <= 16'h0106;    16'd64837: out <= 16'h06C5;    16'd64838: out <= 16'hFFEC;    16'd64839: out <= 16'h0245;
    16'd64840: out <= 16'h04FE;    16'd64841: out <= 16'h0699;    16'd64842: out <= 16'h0333;    16'd64843: out <= 16'h024E;
    16'd64844: out <= 16'h048C;    16'd64845: out <= 16'h0028;    16'd64846: out <= 16'h09ED;    16'd64847: out <= 16'h0077;
    16'd64848: out <= 16'hFF46;    16'd64849: out <= 16'h0384;    16'd64850: out <= 16'h053E;    16'd64851: out <= 16'hFE02;
    16'd64852: out <= 16'h02C4;    16'd64853: out <= 16'h00C2;    16'd64854: out <= 16'h0348;    16'd64855: out <= 16'h0BBA;
    16'd64856: out <= 16'h000E;    16'd64857: out <= 16'h02AC;    16'd64858: out <= 16'h0152;    16'd64859: out <= 16'h02FD;
    16'd64860: out <= 16'hFF21;    16'd64861: out <= 16'h01A1;    16'd64862: out <= 16'h0605;    16'd64863: out <= 16'hFC61;
    16'd64864: out <= 16'hFE95;    16'd64865: out <= 16'h03E5;    16'd64866: out <= 16'hFAC1;    16'd64867: out <= 16'h0A2E;
    16'd64868: out <= 16'h0069;    16'd64869: out <= 16'h019A;    16'd64870: out <= 16'h0063;    16'd64871: out <= 16'hFCF7;
    16'd64872: out <= 16'hFFA3;    16'd64873: out <= 16'h00CD;    16'd64874: out <= 16'hFCB1;    16'd64875: out <= 16'hFA1F;
    16'd64876: out <= 16'h0269;    16'd64877: out <= 16'hFE98;    16'd64878: out <= 16'hF76E;    16'd64879: out <= 16'hFFD7;
    16'd64880: out <= 16'h0604;    16'd64881: out <= 16'hFDA7;    16'd64882: out <= 16'hFFE3;    16'd64883: out <= 16'h0187;
    16'd64884: out <= 16'hFD03;    16'd64885: out <= 16'hFDCE;    16'd64886: out <= 16'hFC5B;    16'd64887: out <= 16'hFF7E;
    16'd64888: out <= 16'h01CA;    16'd64889: out <= 16'h01FA;    16'd64890: out <= 16'h023F;    16'd64891: out <= 16'h0001;
    16'd64892: out <= 16'hFE9B;    16'd64893: out <= 16'hFA63;    16'd64894: out <= 16'hFDDF;    16'd64895: out <= 16'h0198;
    16'd64896: out <= 16'hFF20;    16'd64897: out <= 16'h045C;    16'd64898: out <= 16'hFEFC;    16'd64899: out <= 16'hFB64;
    16'd64900: out <= 16'h0066;    16'd64901: out <= 16'hFC54;    16'd64902: out <= 16'hFFB9;    16'd64903: out <= 16'hFEFE;
    16'd64904: out <= 16'hFDD4;    16'd64905: out <= 16'hFDF5;    16'd64906: out <= 16'hFF6E;    16'd64907: out <= 16'hFFE4;
    16'd64908: out <= 16'h0028;    16'd64909: out <= 16'h03F7;    16'd64910: out <= 16'hF61F;    16'd64911: out <= 16'h01C3;
    16'd64912: out <= 16'hFF74;    16'd64913: out <= 16'hF872;    16'd64914: out <= 16'h01D1;    16'd64915: out <= 16'h01AE;
    16'd64916: out <= 16'h02AC;    16'd64917: out <= 16'hFFC0;    16'd64918: out <= 16'h0142;    16'd64919: out <= 16'hFC9C;
    16'd64920: out <= 16'hFE31;    16'd64921: out <= 16'h0215;    16'd64922: out <= 16'h0085;    16'd64923: out <= 16'hFEE7;
    16'd64924: out <= 16'hFA6B;    16'd64925: out <= 16'h0929;    16'd64926: out <= 16'h0989;    16'd64927: out <= 16'h06D1;
    16'd64928: out <= 16'h03FC;    16'd64929: out <= 16'h0B5F;    16'd64930: out <= 16'h06F8;    16'd64931: out <= 16'h0502;
    16'd64932: out <= 16'h0A1A;    16'd64933: out <= 16'hFB96;    16'd64934: out <= 16'h0BAF;    16'd64935: out <= 16'h09B1;
    16'd64936: out <= 16'h09C2;    16'd64937: out <= 16'h05C5;    16'd64938: out <= 16'h04EF;    16'd64939: out <= 16'hFD2A;
    16'd64940: out <= 16'h0143;    16'd64941: out <= 16'h0CA6;    16'd64942: out <= 16'h01CB;    16'd64943: out <= 16'h0321;
    16'd64944: out <= 16'h08CC;    16'd64945: out <= 16'h01E8;    16'd64946: out <= 16'h05D3;    16'd64947: out <= 16'h0538;
    16'd64948: out <= 16'h057C;    16'd64949: out <= 16'h0060;    16'd64950: out <= 16'h02E6;    16'd64951: out <= 16'h041A;
    16'd64952: out <= 16'h0B3E;    16'd64953: out <= 16'h09A9;    16'd64954: out <= 16'h004C;    16'd64955: out <= 16'hFAA7;
    16'd64956: out <= 16'h046D;    16'd64957: out <= 16'hFDCB;    16'd64958: out <= 16'h043A;    16'd64959: out <= 16'h02B0;
    16'd64960: out <= 16'h0CA3;    16'd64961: out <= 16'h05A7;    16'd64962: out <= 16'h0614;    16'd64963: out <= 16'h03FB;
    16'd64964: out <= 16'h064B;    16'd64965: out <= 16'hFB6D;    16'd64966: out <= 16'hFF61;    16'd64967: out <= 16'h001F;
    16'd64968: out <= 16'hFCC1;    16'd64969: out <= 16'hFA2C;    16'd64970: out <= 16'hFFDB;    16'd64971: out <= 16'h000A;
    16'd64972: out <= 16'h0263;    16'd64973: out <= 16'h0681;    16'd64974: out <= 16'hFE44;    16'd64975: out <= 16'hFBB2;
    16'd64976: out <= 16'hFEC0;    16'd64977: out <= 16'hFC9B;    16'd64978: out <= 16'hFF88;    16'd64979: out <= 16'h0733;
    16'd64980: out <= 16'hFDD5;    16'd64981: out <= 16'hFE84;    16'd64982: out <= 16'h0231;    16'd64983: out <= 16'h0550;
    16'd64984: out <= 16'hFBAF;    16'd64985: out <= 16'h01B3;    16'd64986: out <= 16'hFE60;    16'd64987: out <= 16'h01C8;
    16'd64988: out <= 16'h0245;    16'd64989: out <= 16'h0400;    16'd64990: out <= 16'h0367;    16'd64991: out <= 16'h0132;
    16'd64992: out <= 16'h0004;    16'd64993: out <= 16'hFECE;    16'd64994: out <= 16'hFE30;    16'd64995: out <= 16'h0295;
    16'd64996: out <= 16'hFD86;    16'd64997: out <= 16'h041A;    16'd64998: out <= 16'h038E;    16'd64999: out <= 16'hFCB0;
    16'd65000: out <= 16'h035F;    16'd65001: out <= 16'hFA11;    16'd65002: out <= 16'hFCD7;    16'd65003: out <= 16'hFF95;
    16'd65004: out <= 16'hF937;    16'd65005: out <= 16'hFD06;    16'd65006: out <= 16'hFBEB;    16'd65007: out <= 16'h006D;
    16'd65008: out <= 16'h0111;    16'd65009: out <= 16'hFCAE;    16'd65010: out <= 16'hFD9D;    16'd65011: out <= 16'hF82F;
    16'd65012: out <= 16'h0309;    16'd65013: out <= 16'h031E;    16'd65014: out <= 16'hFF17;    16'd65015: out <= 16'hFF21;
    16'd65016: out <= 16'hFE23;    16'd65017: out <= 16'h0768;    16'd65018: out <= 16'hFEF3;    16'd65019: out <= 16'h01BD;
    16'd65020: out <= 16'h0557;    16'd65021: out <= 16'hFD2D;    16'd65022: out <= 16'h005E;    16'd65023: out <= 16'h003E;
    16'd65024: out <= 16'h03E3;    16'd65025: out <= 16'hFD69;    16'd65026: out <= 16'hFD98;    16'd65027: out <= 16'hFC5F;
    16'd65028: out <= 16'h02D5;    16'd65029: out <= 16'h0380;    16'd65030: out <= 16'hFF7E;    16'd65031: out <= 16'h0053;
    16'd65032: out <= 16'hF7D9;    16'd65033: out <= 16'hF947;    16'd65034: out <= 16'hFEB9;    16'd65035: out <= 16'hFA72;
    16'd65036: out <= 16'h02C9;    16'd65037: out <= 16'h0008;    16'd65038: out <= 16'h0353;    16'd65039: out <= 16'hFD7D;
    16'd65040: out <= 16'h0468;    16'd65041: out <= 16'hFFE0;    16'd65042: out <= 16'h0443;    16'd65043: out <= 16'hFEF3;
    16'd65044: out <= 16'hFED0;    16'd65045: out <= 16'hF855;    16'd65046: out <= 16'hFE1A;    16'd65047: out <= 16'h0528;
    16'd65048: out <= 16'hFD57;    16'd65049: out <= 16'h0483;    16'd65050: out <= 16'h0748;    16'd65051: out <= 16'hFE22;
    16'd65052: out <= 16'h02B4;    16'd65053: out <= 16'hFE76;    16'd65054: out <= 16'h0228;    16'd65055: out <= 16'hFB57;
    16'd65056: out <= 16'h08FA;    16'd65057: out <= 16'hFD16;    16'd65058: out <= 16'h047C;    16'd65059: out <= 16'h03AF;
    16'd65060: out <= 16'h09ED;    16'd65061: out <= 16'h013D;    16'd65062: out <= 16'h02A5;    16'd65063: out <= 16'hFE81;
    16'd65064: out <= 16'h0800;    16'd65065: out <= 16'h0880;    16'd65066: out <= 16'h087E;    16'd65067: out <= 16'h0647;
    16'd65068: out <= 16'h03D6;    16'd65069: out <= 16'h0206;    16'd65070: out <= 16'h002F;    16'd65071: out <= 16'hFD4D;
    16'd65072: out <= 16'h0203;    16'd65073: out <= 16'hFF37;    16'd65074: out <= 16'h0290;    16'd65075: out <= 16'h064A;
    16'd65076: out <= 16'h0ADD;    16'd65077: out <= 16'hFC6C;    16'd65078: out <= 16'h0031;    16'd65079: out <= 16'h0487;
    16'd65080: out <= 16'hFA12;    16'd65081: out <= 16'h0BB3;    16'd65082: out <= 16'h044B;    16'd65083: out <= 16'h06FB;
    16'd65084: out <= 16'h06F4;    16'd65085: out <= 16'h0021;    16'd65086: out <= 16'hFD80;    16'd65087: out <= 16'h0AA5;
    16'd65088: out <= 16'h03C3;    16'd65089: out <= 16'h090A;    16'd65090: out <= 16'h0144;    16'd65091: out <= 16'h03AB;
    16'd65092: out <= 16'h01DB;    16'd65093: out <= 16'h05C2;    16'd65094: out <= 16'h0283;    16'd65095: out <= 16'hFF00;
    16'd65096: out <= 16'h0658;    16'd65097: out <= 16'h0BCC;    16'd65098: out <= 16'h0253;    16'd65099: out <= 16'h08DA;
    16'd65100: out <= 16'h079B;    16'd65101: out <= 16'h0597;    16'd65102: out <= 16'h0007;    16'd65103: out <= 16'h080A;
    16'd65104: out <= 16'h09CE;    16'd65105: out <= 16'h0465;    16'd65106: out <= 16'hFD57;    16'd65107: out <= 16'h033B;
    16'd65108: out <= 16'hFF6B;    16'd65109: out <= 16'h065E;    16'd65110: out <= 16'hFEB4;    16'd65111: out <= 16'h053E;
    16'd65112: out <= 16'h064F;    16'd65113: out <= 16'h07A9;    16'd65114: out <= 16'h06E2;    16'd65115: out <= 16'h0CE2;
    16'd65116: out <= 16'h0640;    16'd65117: out <= 16'h0092;    16'd65118: out <= 16'h06B2;    16'd65119: out <= 16'hFFFE;
    16'd65120: out <= 16'hFAC5;    16'd65121: out <= 16'h0232;    16'd65122: out <= 16'h0053;    16'd65123: out <= 16'hFB99;
    16'd65124: out <= 16'hFAB1;    16'd65125: out <= 16'h0047;    16'd65126: out <= 16'hFD36;    16'd65127: out <= 16'h00F0;
    16'd65128: out <= 16'h0355;    16'd65129: out <= 16'hFFF3;    16'd65130: out <= 16'hFD15;    16'd65131: out <= 16'hFE4F;
    16'd65132: out <= 16'hFD73;    16'd65133: out <= 16'hFEC4;    16'd65134: out <= 16'hFFF8;    16'd65135: out <= 16'hFF0E;
    16'd65136: out <= 16'h00D0;    16'd65137: out <= 16'hFF3E;    16'd65138: out <= 16'hF581;    16'd65139: out <= 16'hFCF2;
    16'd65140: out <= 16'hFEFC;    16'd65141: out <= 16'h0160;    16'd65142: out <= 16'hFF04;    16'd65143: out <= 16'h0730;
    16'd65144: out <= 16'hFD35;    16'd65145: out <= 16'h0376;    16'd65146: out <= 16'h054F;    16'd65147: out <= 16'hFB79;
    16'd65148: out <= 16'hFFBB;    16'd65149: out <= 16'hFD71;    16'd65150: out <= 16'hFCDE;    16'd65151: out <= 16'h0176;
    16'd65152: out <= 16'h0068;    16'd65153: out <= 16'hFC65;    16'd65154: out <= 16'hFF70;    16'd65155: out <= 16'h0752;
    16'd65156: out <= 16'hF582;    16'd65157: out <= 16'hF9F0;    16'd65158: out <= 16'h0780;    16'd65159: out <= 16'h02E4;
    16'd65160: out <= 16'h023A;    16'd65161: out <= 16'h00AA;    16'd65162: out <= 16'hFED7;    16'd65163: out <= 16'hF806;
    16'd65164: out <= 16'h0A82;    16'd65165: out <= 16'h0042;    16'd65166: out <= 16'hFE57;    16'd65167: out <= 16'hFD98;
    16'd65168: out <= 16'hFEFF;    16'd65169: out <= 16'hFC8B;    16'd65170: out <= 16'hFE83;    16'd65171: out <= 16'h08A2;
    16'd65172: out <= 16'h025A;    16'd65173: out <= 16'hFF90;    16'd65174: out <= 16'h017C;    16'd65175: out <= 16'hFF7F;
    16'd65176: out <= 16'hFFEC;    16'd65177: out <= 16'h0148;    16'd65178: out <= 16'h02DC;    16'd65179: out <= 16'h05C9;
    16'd65180: out <= 16'hF9E3;    16'd65181: out <= 16'h063F;    16'd65182: out <= 16'h005A;    16'd65183: out <= 16'h09BF;
    16'd65184: out <= 16'h0753;    16'd65185: out <= 16'hFA6E;    16'd65186: out <= 16'h00BC;    16'd65187: out <= 16'hFFD4;
    16'd65188: out <= 16'h017D;    16'd65189: out <= 16'h0580;    16'd65190: out <= 16'h00C2;    16'd65191: out <= 16'h02FE;
    16'd65192: out <= 16'h045B;    16'd65193: out <= 16'h04C7;    16'd65194: out <= 16'h063A;    16'd65195: out <= 16'h056A;
    16'd65196: out <= 16'h0035;    16'd65197: out <= 16'h0423;    16'd65198: out <= 16'hFF6C;    16'd65199: out <= 16'h01D0;
    16'd65200: out <= 16'h080E;    16'd65201: out <= 16'h03C3;    16'd65202: out <= 16'h0874;    16'd65203: out <= 16'h0853;
    16'd65204: out <= 16'h00BD;    16'd65205: out <= 16'h092D;    16'd65206: out <= 16'h0B3F;    16'd65207: out <= 16'h0471;
    16'd65208: out <= 16'hFE68;    16'd65209: out <= 16'h0D92;    16'd65210: out <= 16'h001A;    16'd65211: out <= 16'h0435;
    16'd65212: out <= 16'h01FD;    16'd65213: out <= 16'h0477;    16'd65214: out <= 16'h017F;    16'd65215: out <= 16'h02C4;
    16'd65216: out <= 16'h0B99;    16'd65217: out <= 16'h082A;    16'd65218: out <= 16'h0ACC;    16'd65219: out <= 16'h05A8;
    16'd65220: out <= 16'hFDC7;    16'd65221: out <= 16'h0407;    16'd65222: out <= 16'hFE80;    16'd65223: out <= 16'h039F;
    16'd65224: out <= 16'h003F;    16'd65225: out <= 16'h026C;    16'd65226: out <= 16'h02C0;    16'd65227: out <= 16'hFB6E;
    16'd65228: out <= 16'h0AEF;    16'd65229: out <= 16'hFD98;    16'd65230: out <= 16'hFCD8;    16'd65231: out <= 16'hF882;
    16'd65232: out <= 16'hFFD2;    16'd65233: out <= 16'hFF6F;    16'd65234: out <= 16'h02A5;    16'd65235: out <= 16'h003D;
    16'd65236: out <= 16'hFE21;    16'd65237: out <= 16'hFA3D;    16'd65238: out <= 16'h00C0;    16'd65239: out <= 16'h0442;
    16'd65240: out <= 16'h0030;    16'd65241: out <= 16'h0777;    16'd65242: out <= 16'h022A;    16'd65243: out <= 16'h01F0;
    16'd65244: out <= 16'hFB67;    16'd65245: out <= 16'h01F1;    16'd65246: out <= 16'h0409;    16'd65247: out <= 16'h03FA;
    16'd65248: out <= 16'hFB2D;    16'd65249: out <= 16'h0508;    16'd65250: out <= 16'hFCC4;    16'd65251: out <= 16'hF93F;
    16'd65252: out <= 16'h009D;    16'd65253: out <= 16'hFA1C;    16'd65254: out <= 16'hF6B7;    16'd65255: out <= 16'h00B1;
    16'd65256: out <= 16'hFDF4;    16'd65257: out <= 16'h01CA;    16'd65258: out <= 16'h0008;    16'd65259: out <= 16'hFFF1;
    16'd65260: out <= 16'h004D;    16'd65261: out <= 16'h04DE;    16'd65262: out <= 16'hFB71;    16'd65263: out <= 16'h0195;
    16'd65264: out <= 16'hFF87;    16'd65265: out <= 16'hFB85;    16'd65266: out <= 16'h0244;    16'd65267: out <= 16'hFFCB;
    16'd65268: out <= 16'h09E7;    16'd65269: out <= 16'hFED6;    16'd65270: out <= 16'hFD46;    16'd65271: out <= 16'h021D;
    16'd65272: out <= 16'hFF29;    16'd65273: out <= 16'h054E;    16'd65274: out <= 16'hFAAC;    16'd65275: out <= 16'hFDBD;
    16'd65276: out <= 16'hFF11;    16'd65277: out <= 16'h017A;    16'd65278: out <= 16'h04E6;    16'd65279: out <= 16'h000D;
    16'd65280: out <= 16'h0065;    16'd65281: out <= 16'h038C;    16'd65282: out <= 16'h0254;    16'd65283: out <= 16'hFCCB;
    16'd65284: out <= 16'h0802;    16'd65285: out <= 16'hFF18;    16'd65286: out <= 16'hFA04;    16'd65287: out <= 16'hFFD3;
    16'd65288: out <= 16'hF327;    16'd65289: out <= 16'hFD9F;    16'd65290: out <= 16'hFEE6;    16'd65291: out <= 16'h0355;
    16'd65292: out <= 16'hFDDA;    16'd65293: out <= 16'hFFDC;    16'd65294: out <= 16'h0128;    16'd65295: out <= 16'h0031;
    16'd65296: out <= 16'h024E;    16'd65297: out <= 16'h0375;    16'd65298: out <= 16'h0433;    16'd65299: out <= 16'hF935;
    16'd65300: out <= 16'hFEA7;    16'd65301: out <= 16'h05B2;    16'd65302: out <= 16'h0296;    16'd65303: out <= 16'hFE63;
    16'd65304: out <= 16'h04C9;    16'd65305: out <= 16'hFC4C;    16'd65306: out <= 16'h03ED;    16'd65307: out <= 16'h0027;
    16'd65308: out <= 16'h005B;    16'd65309: out <= 16'hFDE6;    16'd65310: out <= 16'hFC5B;    16'd65311: out <= 16'h0729;
    16'd65312: out <= 16'h0C4C;    16'd65313: out <= 16'hFA69;    16'd65314: out <= 16'h04B8;    16'd65315: out <= 16'h01E6;
    16'd65316: out <= 16'h08E6;    16'd65317: out <= 16'h08BB;    16'd65318: out <= 16'h0527;    16'd65319: out <= 16'h041A;
    16'd65320: out <= 16'h06DF;    16'd65321: out <= 16'hFD6C;    16'd65322: out <= 16'hFD6F;    16'd65323: out <= 16'hFC51;
    16'd65324: out <= 16'h0607;    16'd65325: out <= 16'h0C53;    16'd65326: out <= 16'h070B;    16'd65327: out <= 16'h0299;
    16'd65328: out <= 16'h0557;    16'd65329: out <= 16'h0998;    16'd65330: out <= 16'h0025;    16'd65331: out <= 16'h07A1;
    16'd65332: out <= 16'h06F3;    16'd65333: out <= 16'h0032;    16'd65334: out <= 16'h0128;    16'd65335: out <= 16'h0210;
    16'd65336: out <= 16'h052C;    16'd65337: out <= 16'h0379;    16'd65338: out <= 16'h0833;    16'd65339: out <= 16'h0854;
    16'd65340: out <= 16'hFEEB;    16'd65341: out <= 16'h02DB;    16'd65342: out <= 16'h0882;    16'd65343: out <= 16'h0274;
    16'd65344: out <= 16'hFD68;    16'd65345: out <= 16'h01A7;    16'd65346: out <= 16'hFE49;    16'd65347: out <= 16'h00F2;
    16'd65348: out <= 16'h0897;    16'd65349: out <= 16'h020A;    16'd65350: out <= 16'h0258;    16'd65351: out <= 16'h07BB;
    16'd65352: out <= 16'h02EC;    16'd65353: out <= 16'h03D7;    16'd65354: out <= 16'h05D0;    16'd65355: out <= 16'h0587;
    16'd65356: out <= 16'h0360;    16'd65357: out <= 16'h04C1;    16'd65358: out <= 16'h09FF;    16'd65359: out <= 16'h02F9;
    16'd65360: out <= 16'h028A;    16'd65361: out <= 16'h020A;    16'd65362: out <= 16'h019D;    16'd65363: out <= 16'hFA8D;
    16'd65364: out <= 16'h0256;    16'd65365: out <= 16'hF8E5;    16'd65366: out <= 16'hFD1B;    16'd65367: out <= 16'h016F;
    16'd65368: out <= 16'hFCF6;    16'd65369: out <= 16'h05BA;    16'd65370: out <= 16'h03D3;    16'd65371: out <= 16'h039E;
    16'd65372: out <= 16'hFFFE;    16'd65373: out <= 16'h01E3;    16'd65374: out <= 16'hFD69;    16'd65375: out <= 16'h0301;
    16'd65376: out <= 16'h0093;    16'd65377: out <= 16'hFF4B;    16'd65378: out <= 16'h04F2;    16'd65379: out <= 16'h01AA;
    16'd65380: out <= 16'h01D1;    16'd65381: out <= 16'h0009;    16'd65382: out <= 16'hFF9C;    16'd65383: out <= 16'h0319;
    16'd65384: out <= 16'h0156;    16'd65385: out <= 16'h05EF;    16'd65386: out <= 16'hF988;    16'd65387: out <= 16'h00E3;
    16'd65388: out <= 16'h0545;    16'd65389: out <= 16'h0518;    16'd65390: out <= 16'hFB73;    16'd65391: out <= 16'h001B;
    16'd65392: out <= 16'hFC04;    16'd65393: out <= 16'hFFC5;    16'd65394: out <= 16'h009F;    16'd65395: out <= 16'hFA42;
    16'd65396: out <= 16'h080F;    16'd65397: out <= 16'h02A8;    16'd65398: out <= 16'hFC87;    16'd65399: out <= 16'hF94A;
    16'd65400: out <= 16'h0325;    16'd65401: out <= 16'hFF04;    16'd65402: out <= 16'hFC9A;    16'd65403: out <= 16'h020B;
    16'd65404: out <= 16'hFB9E;    16'd65405: out <= 16'hFED8;    16'd65406: out <= 16'hFBAD;    16'd65407: out <= 16'h0695;
    16'd65408: out <= 16'h03FC;    16'd65409: out <= 16'hF9B7;    16'd65410: out <= 16'h0261;    16'd65411: out <= 16'h011C;
    16'd65412: out <= 16'h030E;    16'd65413: out <= 16'h0391;    16'd65414: out <= 16'hFE3D;    16'd65415: out <= 16'hFCBD;
    16'd65416: out <= 16'h01A1;    16'd65417: out <= 16'hFF8F;    16'd65418: out <= 16'hFF9A;    16'd65419: out <= 16'h0419;
    16'd65420: out <= 16'h03BA;    16'd65421: out <= 16'hFE51;    16'd65422: out <= 16'hFC73;    16'd65423: out <= 16'hFDD9;
    16'd65424: out <= 16'h0186;    16'd65425: out <= 16'h0707;    16'd65426: out <= 16'hFB55;    16'd65427: out <= 16'h0137;
    16'd65428: out <= 16'h009A;    16'd65429: out <= 16'h03C2;    16'd65430: out <= 16'h0275;    16'd65431: out <= 16'hFF40;
    16'd65432: out <= 16'h01EC;    16'd65433: out <= 16'hFD96;    16'd65434: out <= 16'hFF29;    16'd65435: out <= 16'hFCBA;
    16'd65436: out <= 16'h07B8;    16'd65437: out <= 16'hFFA2;    16'd65438: out <= 16'hFF29;    16'd65439: out <= 16'h0466;
    16'd65440: out <= 16'h06EA;    16'd65441: out <= 16'h02F9;    16'd65442: out <= 16'h0CB4;    16'd65443: out <= 16'h0617;
    16'd65444: out <= 16'h044C;    16'd65445: out <= 16'h0676;    16'd65446: out <= 16'h0772;    16'd65447: out <= 16'h05F9;
    16'd65448: out <= 16'hFF12;    16'd65449: out <= 16'h0282;    16'd65450: out <= 16'h0A37;    16'd65451: out <= 16'h049E;
    16'd65452: out <= 16'h08D5;    16'd65453: out <= 16'h00A5;    16'd65454: out <= 16'h0303;    16'd65455: out <= 16'h0263;
    16'd65456: out <= 16'hFEB7;    16'd65457: out <= 16'h01E3;    16'd65458: out <= 16'h03F7;    16'd65459: out <= 16'h0503;
    16'd65460: out <= 16'h05A2;    16'd65461: out <= 16'h0568;    16'd65462: out <= 16'hFDFC;    16'd65463: out <= 16'h04CD;
    16'd65464: out <= 16'h09CC;    16'd65465: out <= 16'h0C1B;    16'd65466: out <= 16'h0084;    16'd65467: out <= 16'h0182;
    16'd65468: out <= 16'h069C;    16'd65469: out <= 16'h0977;    16'd65470: out <= 16'h0019;    16'd65471: out <= 16'h0250;
    16'd65472: out <= 16'h0234;    16'd65473: out <= 16'h0476;    16'd65474: out <= 16'hFFDE;    16'd65475: out <= 16'h0C63;
    16'd65476: out <= 16'h09C6;    16'd65477: out <= 16'hFF7A;    16'd65478: out <= 16'hFDEB;    16'd65479: out <= 16'hFA2C;
    16'd65480: out <= 16'h0039;    16'd65481: out <= 16'h078C;    16'd65482: out <= 16'hFFDC;    16'd65483: out <= 16'hFB00;
    16'd65484: out <= 16'hFAE1;    16'd65485: out <= 16'hFE05;    16'd65486: out <= 16'h01AA;    16'd65487: out <= 16'hFCF3;
    16'd65488: out <= 16'h056C;    16'd65489: out <= 16'h005B;    16'd65490: out <= 16'hFAA5;    16'd65491: out <= 16'h03C0;
    16'd65492: out <= 16'h032E;    16'd65493: out <= 16'hFC23;    16'd65494: out <= 16'h0079;    16'd65495: out <= 16'hFEBA;
    16'd65496: out <= 16'h0057;    16'd65497: out <= 16'hFCD9;    16'd65498: out <= 16'h02A9;    16'd65499: out <= 16'h0555;
    16'd65500: out <= 16'h04BC;    16'd65501: out <= 16'h01C2;    16'd65502: out <= 16'hFA09;    16'd65503: out <= 16'h03C2;
    16'd65504: out <= 16'h00B8;    16'd65505: out <= 16'hFE07;    16'd65506: out <= 16'hFCC3;    16'd65507: out <= 16'h0119;
    16'd65508: out <= 16'h032F;    16'd65509: out <= 16'hFF4B;    16'd65510: out <= 16'h02BC;    16'd65511: out <= 16'hFD56;
    16'd65512: out <= 16'hFA2E;    16'd65513: out <= 16'hFFE4;    16'd65514: out <= 16'h0004;    16'd65515: out <= 16'h01FF;
    16'd65516: out <= 16'hF821;    16'd65517: out <= 16'h0044;    16'd65518: out <= 16'hFFDB;    16'd65519: out <= 16'h032B;
    16'd65520: out <= 16'hFBD2;    16'd65521: out <= 16'hF836;    16'd65522: out <= 16'h04D7;    16'd65523: out <= 16'hFBA1;
    16'd65524: out <= 16'hF93A;    16'd65525: out <= 16'h0866;    16'd65526: out <= 16'h0182;    16'd65527: out <= 16'h000A;
    16'd65528: out <= 16'hFE76;    16'd65529: out <= 16'hFE1F;    16'd65530: out <= 16'h0162;    16'd65531: out <= 16'h025E;
    16'd65532: out <= 16'hFE47;    16'd65533: out <= 16'hFA6C;    16'd65534: out <= 16'hFD2A;    16'd65535: out <= 16'hF7E9;
    default: out <= 16'h0000;
    endcase
endmodule
